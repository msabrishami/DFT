1 N1 0 5 0
1 N5 0 5 0
1 N9 0 6 0
1 N13 0 6 0
1 N17 0 6 0
1 N21 0 6 0
1 N25 0 6 0
1 N29 0 4 0
1 N33 0 6 0
1 N37 0 6 0
1 N41 0 5 0
1 N45 0 4 0
1 N49 0 6 0
1 N53 0 5 0
1 N57 0 6 0
1 N61 0 6 0
1 N65 0 5 0
1 N69 0 6 0
1 N73 0 6 0
1 N77 0 5 0
1 N81 0 6 0
1 N85 0 6 0
1 N89 0 5 0
1 N93 0 5 0
1 N97 0 6 0
1 N101 0 5 0
1 N105 0 6 0
1 N109 0 5 0
1 N113 0 6 0
1 N117 0 5 0
1 N121 0 6 0
1 N125 0 5 0
1 N129 0 1 0
1 N130 0 1 0
1 N131 0 1 0
1 N132 0 1 0
1 N133 0 1 0
1 N134 0 1 0
1 N135 0 1 0
1 N136 0 1 0
1 N137 0 8 0
2 N1-1 1 N1 
2 N1-2 1 N1 
2 N1-3 1 N1 
2 N1-4 1 N1 
2 N1-5 1 N1 
2 N5-1 1 N5 
2 N5-2 1 N5 
2 N5-3 1 N5 
2 N5-4 1 N5 
2 N5-5 1 N5 
2 N9-1 1 N9 
2 N9-2 1 N9 
2 N9-3 1 N9 
2 N9-4 1 N9 
2 N9-5 1 N9 
2 N9-6 1 N9 
2 N13-1 1 N13 
2 N13-2 1 N13 
2 N13-3 1 N13 
2 N13-4 1 N13 
2 N13-5 1 N13 
2 N13-6 1 N13 
2 N17-1 1 N17 
2 N17-2 1 N17 
2 N17-3 1 N17 
2 N17-4 1 N17 
2 N17-5 1 N17 
2 N17-6 1 N17 
2 N21-1 1 N21 
2 N21-2 1 N21 
2 N21-3 1 N21 
2 N21-4 1 N21 
2 N21-5 1 N21 
2 N21-6 1 N21 
2 N25-1 1 N25 
2 N25-2 1 N25 
2 N25-3 1 N25 
2 N25-4 1 N25 
2 N25-5 1 N25 
2 N25-6 1 N25 
2 N29-1 1 N29 
2 N29-2 1 N29 
2 N29-3 1 N29 
2 N29-4 1 N29 
2 N33-1 1 N33 
2 N33-2 1 N33 
2 N33-3 1 N33 
2 N33-4 1 N33 
2 N33-5 1 N33 
2 N33-6 1 N33 
2 N37-1 1 N37 
2 N37-2 1 N37 
2 N37-3 1 N37 
2 N37-4 1 N37 
2 N37-5 1 N37 
2 N37-6 1 N37 
2 N41-1 1 N41 
2 N41-2 1 N41 
2 N41-3 1 N41 
2 N41-4 1 N41 
2 N41-5 1 N41 
2 N45-1 1 N45 
2 N45-2 1 N45 
2 N45-3 1 N45 
2 N45-4 1 N45 
2 N49-1 1 N49 
2 N49-2 1 N49 
2 N49-3 1 N49 
2 N49-4 1 N49 
2 N49-5 1 N49 
2 N49-6 1 N49 
2 N53-1 1 N53 
2 N53-2 1 N53 
2 N53-3 1 N53 
2 N53-4 1 N53 
2 N53-5 1 N53 
2 N57-1 1 N57 
2 N57-2 1 N57 
2 N57-3 1 N57 
2 N57-4 1 N57 
2 N57-5 1 N57 
2 N57-6 1 N57 
2 N61-1 1 N61 
2 N61-2 1 N61 
2 N61-3 1 N61 
2 N61-4 1 N61 
2 N61-5 1 N61 
2 N61-6 1 N61 
2 N65-1 1 N65 
2 N65-2 1 N65 
2 N65-3 1 N65 
2 N65-4 1 N65 
2 N65-5 1 N65 
2 N69-1 1 N69 
2 N69-2 1 N69 
2 N69-3 1 N69 
2 N69-4 1 N69 
2 N69-5 1 N69 
2 N69-6 1 N69 
2 N73-1 1 N73 
2 N73-2 1 N73 
2 N73-3 1 N73 
2 N73-4 1 N73 
2 N73-5 1 N73 
2 N73-6 1 N73 
2 N77-1 1 N77 
2 N77-2 1 N77 
2 N77-3 1 N77 
2 N77-4 1 N77 
2 N77-5 1 N77 
2 N81-1 1 N81 
2 N81-2 1 N81 
2 N81-3 1 N81 
2 N81-4 1 N81 
2 N81-5 1 N81 
2 N81-6 1 N81 
2 N85-1 1 N85 
2 N85-2 1 N85 
2 N85-3 1 N85 
2 N85-4 1 N85 
2 N85-5 1 N85 
2 N85-6 1 N85 
2 N89-1 1 N89 
2 N89-2 1 N89 
2 N89-3 1 N89 
2 N89-4 1 N89 
2 N89-5 1 N89 
2 N93-1 1 N93 
2 N93-2 1 N93 
2 N93-3 1 N93 
2 N93-4 1 N93 
2 N93-5 1 N93 
2 N97-1 1 N97 
2 N97-2 1 N97 
2 N97-3 1 N97 
2 N97-4 1 N97 
2 N97-5 1 N97 
2 N97-6 1 N97 
2 N101-1 1 N101 
2 N101-2 1 N101 
2 N101-3 1 N101 
2 N101-4 1 N101 
2 N101-5 1 N101 
2 N105-1 1 N105 
2 N105-2 1 N105 
2 N105-3 1 N105 
2 N105-4 1 N105 
2 N105-5 1 N105 
2 N105-6 1 N105 
2 N109-1 1 N109 
2 N109-2 1 N109 
2 N109-3 1 N109 
2 N109-4 1 N109 
2 N109-5 1 N109 
2 N113-1 1 N113 
2 N113-2 1 N113 
2 N113-3 1 N113 
2 N113-4 1 N113 
2 N113-5 1 N113 
2 N113-6 1 N113 
2 N117-1 1 N117 
2 N117-2 1 N117 
2 N117-3 1 N117 
2 N117-4 1 N117 
2 N117-5 1 N117 
2 N121-1 1 N121 
2 N121-2 1 N121 
2 N121-3 1 N121 
2 N121-4 1 N121 
2 N121-5 1 N121 
2 N121-6 1 N121 
2 N125-1 1 N125 
2 N125-2 1 N125 
2 N125-3 1 N125 
2 N125-4 1 N125 
2 N125-5 1 N125 
2 N137-1 1 N137 
2 N137-2 1 N137 
2 N137-3 1 N137 
2 N137-4 1 N137 
2 N137-5 1 N137 
2 N137-6 1 N137 
2 N137-7 1 N137 
2 N137-8 1 N137 
0 n595 6 2 2 N129 N137-1
0 n628 6 3 2 N131 N137-2
0 n674 6 3 2 N132 N137-3
0 n719 6 3 2 N130 N137-4
0 n782 6 2 2 N135 N137-5
0 n745 5 3 1 N121-5
0 n599 5 2 1 N89-5
0 n653 5 3 1 N105-5
0 n640 5 3 1 N73-6
0 n793 5 2 1 N5-4
0 n639 5 2 1 N65-5
0 n697 5 3 1 N113-5
0 n650 5 3 1 N97-6
0 n763 5 4 1 N1-5
0 n694 5 3 1 N81-6
0 n693 5 3 1 N13-5
0 n649 5 3 1 N9-6
0 n809 6 2 2 N133 N137-6
0 n779 5 3 1 N45-4
0 n579 5 3 1 N85-6
0 n853 6 2 2 N134 N137-7
0 n758 5 3 1 N33-5
0 n721 5 4 1 N101-5
0 n778 5 2 1 N41-4
0 n584 5 3 1 N69-6
0 n698 5 4 1 N117-5
0 n740 5 4 1 N125-5
0 n802 5 3 1 N29-3
0 n600 5 2 1 N93-5
0 n741 5 3 1 N21-5
0 n654 5 3 1 N25-6
0 n885 6 3 2 N136 N137-8
0 n744 5 4 1 N109-5
0 n578 5 4 1 N77-5
0 n833 5 3 1 N17-5
0 n859 5 3 1 N49-6
0 n873 5 4 1 N53-4
0 n850 5 3 1 N61-6
2 n595-1 1 n595 
2 n595-2 1 n595 
2 n628-1 1 n628 
2 n628-2 1 n628 
2 n628-3 1 n628 
2 n674-1 1 n674 
2 n674-2 1 n674 
2 n674-3 1 n674 
2 n719-1 1 n719 
2 n719-2 1 n719 
2 n719-3 1 n719 
2 n782-1 1 n782 
2 n782-2 1 n782 
2 n745-1 1 n745 
2 n745-2 1 n745 
2 n745-3 1 n745 
2 n599-1 1 n599 
2 n599-2 1 n599 
2 n653-1 1 n653 
2 n653-2 1 n653 
2 n653-3 1 n653 
2 n640-1 1 n640 
2 n640-2 1 n640 
2 n640-3 1 n640 
2 n793-1 1 n793 
2 n793-2 1 n793 
2 n639-1 1 n639 
2 n639-2 1 n639 
2 n697-1 1 n697 
2 n697-2 1 n697 
2 n697-3 1 n697 
2 n650-1 1 n650 
2 n650-2 1 n650 
2 n650-3 1 n650 
2 n763-1 1 n763 
2 n763-2 1 n763 
2 n763-3 1 n763 
2 n763-4 1 n763 
2 n694-1 1 n694 
2 n694-2 1 n694 
2 n694-3 1 n694 
2 n693-1 1 n693 
2 n693-2 1 n693 
2 n693-3 1 n693 
2 n649-1 1 n649 
2 n649-2 1 n649 
2 n649-3 1 n649 
2 n809-1 1 n809 
2 n809-2 1 n809 
2 n779-1 1 n779 
2 n779-2 1 n779 
2 n779-3 1 n779 
2 n579-1 1 n579 
2 n579-2 1 n579 
2 n579-3 1 n579 
2 n853-1 1 n853 
2 n853-2 1 n853 
2 n758-1 1 n758 
2 n758-2 1 n758 
2 n758-3 1 n758 
2 n721-1 1 n721 
2 n721-2 1 n721 
2 n721-3 1 n721 
2 n721-4 1 n721 
2 n778-1 1 n778 
2 n778-2 1 n778 
2 n584-1 1 n584 
2 n584-2 1 n584 
2 n584-3 1 n584 
2 n698-1 1 n698 
2 n698-2 1 n698 
2 n698-3 1 n698 
2 n698-4 1 n698 
2 n740-1 1 n740 
2 n740-2 1 n740 
2 n740-3 1 n740 
2 n740-4 1 n740 
2 n802-1 1 n802 
2 n802-2 1 n802 
2 n802-3 1 n802 
2 n600-1 1 n600 
2 n600-2 1 n600 
2 n741-1 1 n741 
2 n741-2 1 n741 
2 n741-3 1 n741 
2 n654-1 1 n654 
2 n654-2 1 n654 
2 n654-3 1 n654 
2 n885-1 1 n885 
2 n885-2 1 n885 
2 n885-3 1 n885 
2 n744-1 1 n744 
2 n744-2 1 n744 
2 n744-3 1 n744 
2 n744-4 1 n744 
2 n578-1 1 n578 
2 n578-2 1 n578 
2 n578-3 1 n578 
2 n578-4 1 n578 
2 n833-1 1 n833 
2 n833-2 1 n833 
2 n833-3 1 n833 
2 n859-1 1 n859 
2 n859-2 1 n859 
2 n859-3 1 n859 
2 n873-1 1 n873 
2 n873-2 1 n873 
2 n873-3 1 n873 
2 n873-4 1 n873 
2 n850-1 1 n850 
2 n850-2 1 n850 
2 n850-3 1 n850 
0 n577 6 1 2 N85-3 n578-1
0 n576 6 1 2 N77-3 n579-1
0 n598 6 1 2 N93-3 n599-1
0 n597 6 1 2 N89-3 n600-1
0 n612 4 1 2 N85-4 n578-2
0 n611 4 1 2 N77-4 n579-2
0 n638 6 1 2 N73-3 n639-1
0 n637 6 1 2 N65-3 n640-1
0 n625 5 2 1 n628-2
0 n648 6 1 2 N97-3 n649-1
0 n647 6 1 2 N9-3 n650-1
0 n652 4 1 2 N25-3 n653-1
0 n651 4 1 2 N105-3 n654-1
0 n658 6 1 2 N25-4 n653-2
0 n657 6 1 2 N105-4 n654-2
0 n660 4 1 2 N97-4 n649-2
0 n659 4 1 2 N9-4 n650-2
0 n671 5 2 1 n674-2
0 n692 6 1 2 N81-3 n693-1
0 n691 6 1 2 N13-3 n694-1
0 n696 4 1 2 N117-3 n697-1
0 n695 4 1 2 N113-3 n698-1
0 n702 6 1 2 N117-4 n697-2
0 n701 6 1 2 N113-4 n698-2
0 n704 4 1 2 N81-4 n693-2
0 n703 4 1 2 N13-4 n694-2
0 n718 6 1 2 N101-3 n719-1
0 n733 4 1 2 N101-4 n719-2
0 n720 5 2 1 n719-3
0 n739 6 1 2 N21-3 n740-1
0 n738 6 1 2 N125-3 n741-1
0 n743 4 1 2 N121-3 n744-1
0 n742 4 1 2 N109-3 n745-1
0 n749 6 1 2 N121-4 n744-2
0 n748 6 1 2 N109-4 n745-2
0 n751 4 1 2 N21-4 n740-2
0 n750 4 1 2 N125-4 n741-2
0 n757 6 1 2 N73-4 n758-1
0 n756 6 1 2 N33-3 n640-2
0 n777 6 1 2 N45-3 n778-1
0 n776 6 1 2 N41-3 n779-1
0 n781 6 1 2 N37-3 n782-1
0 n780 3 1 2 N37-4 n782-2
0 n790 6 1 2 N89-4 n745-3
0 n789 6 1 2 N121-6 n599-2
0 n792 6 1 2 N5-3 n653-3
0 n791 6 1 2 N105-6 n793-1
0 n795 4 1 2 N73-5 n758-2
0 n794 4 1 2 N33-4 n640-3
0 n805 6 1 2 N65-4 n793-2
0 n804 6 1 2 N5-5 n639-2
0 n827 6 1 2 N97-5 n697-3
0 n826 6 1 2 N113-6 n650-3
0 n832 6 1 2 N81-5 n833-1
0 n831 6 1 2 N17-3 n694-3
0 n837 6 1 2 N9-5 n693-3
0 n836 6 1 2 N13-6 n649-3
0 n849 6 1 2 N85-5 n850-1
0 n848 6 1 2 N61-3 n579-3
0 n852 6 1 2 N57-3 n853-1
0 n851 3 1 2 N57-4 n853-2
0 n858 6 1 2 N49-3 n758-3
0 n857 6 1 2 N33-6 n859-1
0 n867 6 1 2 N69-5 n778-2
0 n866 6 1 2 N41-5 n584-3
0 n872 3 1 2 N37-5 n873-1
0 n871 6 1 2 N37-6 n873-2
0 n896 6 1 2 N93-4 n802-3
0 n895 6 1 2 N29-4 n600-2
0 n898 6 1 2 N25-5 n741-3
0 n897 6 1 2 N21-6 n654-3
0 n884 5 2 1 n885-2
0 n905 3 1 2 N57-5 n578-3
0 n904 6 1 2 N57-6 n578-4
0 n911 6 1 2 N61-4 n873-3
0 n910 6 1 2 N53-3 n850-2
0 n913 4 1 2 N49-4 n833-2
0 n912 4 1 2 N17-4 n859-2
0 n917 6 1 2 N49-5 n833-3
0 n916 6 1 2 N17-6 n859-3
0 n919 4 1 2 N61-5 n873-4
0 n918 4 1 2 N53-5 n850-3
0 n575 6 1 2 n576 n577
0 n596 6 2 2 n597 n598
0 n585 4 1 2 n611 n612
0 n607 6 4 2 n637 n638
0 n646 6 1 2 n647 n648
0 n645 4 1 2 n651 n652
0 n656 6 1 2 n657 n658
0 n655 4 1 2 n659 n660
0 n690 6 1 2 n691 n692
0 n689 4 1 2 n695 n696
0 n700 6 1 2 n701 n702
0 n699 4 1 2 n703 n704
0 n737 6 1 2 n738 n739
0 n736 4 1 2 n742 n743
0 n747 6 1 2 n748 n749
0 n746 4 1 2 n750 n751
0 n755 6 1 2 n756 n757
0 n774 6 2 2 n776 n777
0 n775 7 2 2 n780 n781
0 n679 6 4 2 n789 n790
0 n724 6 4 2 n791 n792
0 n764 4 1 2 n794 n795
0 n803 6 2 2 n804 n805
0 n726 6 5 2 n826 n827
0 n830 6 2 2 n831 n832
0 n817 6 3 2 n836 n837
0 n847 6 2 2 n848 n849
0 n844 6 2 2 n851 n852
0 n609 6 2 2 n857 n858
0 n865 6 2 2 n866 n867
0 n870 6 2 2 n871 n872
0 n894 6 2 2 n895 n896
0 n816 6 5 2 n897 n898
0 n903 6 2 2 n904 n905
0 n909 6 1 2 n910 n911
0 n908 4 1 2 n912 n913
0 n915 6 1 2 n916 n917
0 n914 4 1 2 n918 n919
2 n625-1 1 n625 
2 n625-2 1 n625 
2 n671-1 1 n671 
2 n671-2 1 n671 
2 n720-1 1 n720 
2 n720-2 1 n720 
2 n884-1 1 n884 
2 n884-2 1 n884 
0 n644 6 1 2 n645 n646
0 n643 6 1 2 n655 n656
0 n688 6 1 2 n689 n690
0 n687 6 1 2 n699 n700
0 n717 6 1 2 n720-1 n721-1
0 n732 4 1 2 n720-2 n721-2
0 n735 6 1 2 n736 n737
0 n734 6 1 2 n746 n747
0 n907 6 1 2 n908 n909
0 n906 6 1 2 n914 n915
2 n596-1 1 n596 
2 n596-2 1 n596 
2 n607-1 1 n607 
2 n607-2 1 n607 
2 n607-3 1 n607 
2 n607-4 1 n607 
2 n774-1 1 n774 
2 n774-2 1 n774 
2 n775-1 1 n775 
2 n775-2 1 n775 
2 n679-1 1 n679 
2 n679-2 1 n679 
2 n679-3 1 n679 
2 n679-4 1 n679 
2 n724-1 1 n724 
2 n724-2 1 n724 
2 n724-3 1 n724 
2 n724-4 1 n724 
2 n803-1 1 n803 
2 n803-2 1 n803 
2 n726-1 1 n726 
2 n726-2 1 n726 
2 n726-3 1 n726 
2 n726-4 1 n726 
2 n726-5 1 n726 
2 n830-1 1 n830 
2 n830-2 1 n830 
2 n817-1 1 n817 
2 n817-2 1 n817 
2 n817-3 1 n817 
2 n847-1 1 n847 
2 n847-2 1 n847 
2 n844-1 1 n844 
2 n844-2 1 n844 
2 n609-1 1 n609 
2 n609-2 1 n609 
2 n865-1 1 n865 
2 n865-2 1 n865 
2 n870-1 1 n870 
2 n870-2 1 n870 
2 n894-1 1 n894 
2 n894-2 1 n894 
2 n816-1 1 n816 
2 n816-2 1 n816 
2 n816-3 1 n816 
2 n816-4 1 n816 
2 n816-5 1 n816 
2 n903-1 1 n903 
2 n903-2 1 n903 
0 n594 3 1 2 n595-1 n596-1
0 n593 6 1 2 n595-2 n596-2
0 n610 5 3 1 n607-3
0 n618 6 2 2 n643 n644
0 n664 6 2 2 n687 n688
0 n716 6 1 2 n717 n718
0 n728 4 1 2 n732 n733
0 n712 6 2 2 n734 n735
0 n773 6 1 2 n774-1 n775-1
0 n772 3 1 2 n774-2 n775-2
0 n727 5 3 1 n724-3
0 n678 5 3 1 n679-4
0 n801 3 1 2 n803-1 n802-1
0 n800 6 1 2 n803-2 n802-2
0 n725 5 4 1 n726-5
0 n829 3 1 2 n763-3 n830-1
0 n828 6 1 2 n763-4 n830-2
0 n785 5 4 1 n817-2
0 n846 3 1 2 n779-2 n847-1
0 n845 6 1 2 n779-3 n847-2
0 n608 5 3 1 n609-2
0 n864 3 1 2 n721-3 n865-1
0 n863 6 1 2 n721-4 n865-2
0 n869 3 1 2 n698-3 n870-1
0 n868 6 1 2 n698-4 n870-2
0 n818 5 4 1 n816-4
0 n893 3 1 2 n740-3 n894-1
0 n892 6 1 2 n740-4 n894-2
0 n902 3 1 2 n744-3 n903-1
0 n901 6 1 2 n744-4 n903-2
0 n877 6 2 2 n906 n907
0 n591 6 2 2 n593 n594
0 n770 6 2 2 n772 n773
0 n798 6 2 2 n800 n801
0 n821 6 3 2 n828 n829
0 n677 6 3 2 n845 n846
0 n631 6 4 2 n863 n864
0 n862 6 2 2 n868 n869
0 n673 6 5 2 n892 n893
0 n627 6 5 2 n901 n902
2 n610-1 1 n610 
2 n610-2 1 n610 
2 n610-3 1 n610 
2 n618-1 1 n618 
2 n618-2 1 n618 
2 n664-1 1 n664 
2 n664-2 1 n664 
2 n712-1 1 n712 
2 n712-2 1 n712 
2 n727-1 1 n727 
2 n727-2 1 n727 
2 n727-3 1 n727 
2 n678-1 1 n678 
2 n678-2 1 n678 
2 n678-3 1 n678 
2 n725-1 1 n725 
2 n725-2 1 n725 
2 n725-3 1 n725 
2 n725-4 1 n725 
2 n785-1 1 n785 
2 n785-2 1 n785 
2 n785-3 1 n785 
2 n785-4 1 n785 
2 n608-1 1 n608 
2 n608-2 1 n608 
2 n608-3 1 n608 
2 n818-1 1 n818 
2 n818-2 1 n818 
2 n818-3 1 n818 
2 n818-4 1 n818 
2 n877-1 1 n877 
2 n877-2 1 n877 
0 n606 6 1 2 n607-1 n608-1
0 n605 6 1 2 n610-1 n609-1
0 n723 4 1 2 n724-1 n725-1
0 n722 4 1 2 n727-1 n726-1
0 n731 6 1 2 n724-2 n725-2
0 n730 6 1 2 n727-2 n726-2
0 n788 6 1 2 n727-3 n679-3
0 n787 6 1 2 n678-3 n724-4
0 n815 6 1 2 n785-3 n816-1
0 n814 6 1 2 n817-1 n818-1
0 n835 4 1 2 n785-4 n816-2
0 n834 4 1 2 n817-3 n818-2
2 n591-1 1 n591 
2 n591-2 1 n591 
2 n770-1 1 n770 
2 n770-2 1 n770 
2 n798-1 1 n798 
2 n798-2 1 n798 
2 n821-1 1 n821 
2 n821-2 1 n821 
2 n821-3 1 n821 
2 n677-1 1 n677 
2 n677-2 1 n677 
2 n677-3 1 n677 
2 n631-1 1 n631 
2 n631-2 1 n631 
2 n631-3 1 n631 
2 n631-4 1 n631 
2 n862-1 1 n862 
2 n862-2 1 n862 
2 n673-1 1 n673 
2 n673-2 1 n673 
2 n673-3 1 n673 
2 n673-4 1 n673 
2 n673-5 1 n673 
2 n627-1 1 n627 
2 n627-2 1 n627 
2 n627-3 1 n627 
2 n627-4 1 n627 
2 n627-5 1 n627 
0 n604 6 2 2 n605 n606
0 n623 6 1 2 n628-1 n627-1
0 n630 4 1 2 n610-2 n631-1
0 n636 6 1 2 n610-3 n631-2
0 n641 4 1 2 n628-3 n627-2
0 n669 6 1 2 n674-1 n673-1
0 n676 4 1 2 n678-1 n677-1
0 n684 6 1 2 n678-2 n677-2
0 n685 4 1 2 n674-3 n673-2
0 n715 4 1 2 n722 n723
0 n729 6 1 2 n730 n731
0 n786 6 2 2 n787 n788
0 n813 6 1 2 n814 n815
0 n819 4 1 2 n725-3 n821-1
0 n603 5 4 1 n821-2
0 n824 6 1 2 n725-4 n821-3
0 n822 4 1 2 n834 n835
0 n680 5 4 1 n677-3
0 n707 5 3 1 n862-1
0 n632 5 3 1 n631-4
0 n882 6 1 2 n885-1 n627-3
0 n887 4 1 2 n818-3 n673-3
0 n891 6 1 2 n818-4 n673-4
0 n672 5 4 1 n673-5
0 n626 5 4 1 n627-4
0 n899 4 1 2 n885-3 n627-5
0 n714 6 1 2 n715 n716
0 n713 6 1 2 n728 n729
2 n604-1 1 n604 
2 n604-2 1 n604 
2 n786-1 1 n786 
2 n786-2 1 n786 
2 n603-1 1 n603 
2 n603-2 1 n603 
2 n603-3 1 n603 
2 n603-4 1 n603 
2 n680-1 1 n680 
2 n680-2 1 n680 
2 n680-3 1 n680 
2 n680-4 1 n680 
2 n707-1 1 n707 
2 n707-2 1 n707 
2 n707-3 1 n707 
2 n632-1 1 n632 
2 n632-2 1 n632 
2 n632-3 1 n632 
2 n672-1 1 n672 
2 n672-2 1 n672 
2 n672-3 1 n672 
2 n672-4 1 n672 
2 n626-1 1 n626 
2 n626-2 1 n626 
2 n626-3 1 n626 
2 n626-4 1 n626 
0 n602 3 1 2 n604-1 n603-1
0 n601 6 1 2 n604-2 n603-2
0 n624 6 1 2 n625-1 n626-1
0 n629 4 1 2 n607-2 n632-1
0 n635 6 1 2 n607-4 n632-2
0 n642 4 1 2 n625-2 n626-2
0 n670 6 1 2 n671-1 n672-1
0 n675 4 1 2 n679-1 n680-1
0 n683 6 1 2 n679-2 n680-2
0 n686 4 1 2 n671-2 n672-2
0 n711 7 2 2 n713 n714
0 n784 3 1 2 n786-1 n785-1
0 n783 6 1 2 n786-2 n785-2
0 n820 4 1 2 n603-3 n726-3
0 n825 6 1 2 n603-4 n726-4
0 n843 3 1 2 n680-3 n844-1
0 n842 6 1 2 n680-4 n844-2
0 n861 6 1 2 n707-3 n631-3
0 n860 6 1 2 n632-3 n862-2
0 n883 6 1 2 n626-3 n884-1
0 n886 4 1 2 n672-3 n816-3
0 n890 6 1 2 n672-4 n816-5
0 n900 4 1 2 n626-4 n884-2
0 n592 7 2 2 n601 n602
0 n622 6 1 2 n623 n624
0 n621 4 1 2 n629 n630
0 n634 6 1 2 n635 n636
0 n633 4 1 2 n641 n642
0 n668 6 1 2 n669 n670
0 n667 4 1 2 n675 n676
0 n682 6 1 2 n683 n684
0 n681 4 1 2 n685 n686
0 n771 7 2 2 n783 n784
0 n812 4 1 2 n819 n820
0 n823 6 1 2 n824 n825
0 n840 6 2 2 n842 n843
0 n856 6 2 2 n860 n861
0 n881 6 1 2 n882 n883
0 n880 4 1 2 n886 n887
0 n889 6 1 2 n890 n891
0 n888 4 1 2 n899 n900
2 n711-1 1 n711 
2 n711-2 1 n711 
0 n620 6 1 2 n621 n622
0 n619 6 1 2 n633 n634
0 n666 6 1 2 n667 n668
0 n665 6 1 2 n681 n682
0 n710 6 1 2 n711-1 n712-1
0 n709 3 1 2 n711-2 n712-2
0 n811 6 1 2 n812 n813
0 n810 6 1 2 n822 n823
0 n879 6 1 2 n880 n881
0 n878 6 1 2 n888 n889
2 n592-1 1 n592 
2 n592-2 1 n592 
2 n771-1 1 n771 
2 n771-2 1 n771 
2 n840-1 1 n840 
2 n840-2 1 n840 
2 n856-1 1 n856 
2 n856-2 1 n856 
0 n590 6 1 2 n591-1 n592-1
0 n589 3 1 2 n591-2 n592-2
0 n617 7 2 2 n619 n620
0 n663 7 2 2 n665 n666
0 n708 6 2 2 n709 n710
0 n769 6 1 2 n770-1 n771-1
0 n768 3 1 2 n770-2 n771-2
0 n808 7 2 2 n810 n811
0 n855 3 1 2 n608-2 n856-1
0 n854 6 1 2 n608-3 n856-2
0 n876 7 2 2 n878 n879
0 n583 6 3 2 n589 n590
0 n762 6 3 2 n768 n769
0 n841 7 2 2 n854 n855
2 n617-1 1 n617 
2 n617-2 1 n617 
2 n663-1 1 n663 
2 n663-2 1 n663 
2 n708-1 1 n708 
2 n708-2 1 n708 
2 n808-1 1 n808 
2 n808-2 1 n808 
2 n876-1 1 n876 
2 n876-2 1 n876 
0 n616 6 1 2 n617-1 n618-1
0 n615 3 1 2 n617-2 n618-2
0 n662 6 1 2 n663-1 n664-1
0 n661 3 1 2 n663-2 n664-2
0 n706 3 1 2 n708-1 n707-1
0 n705 6 1 2 n708-2 n707-2
0 n807 6 1 2 n808-1 n809-1
0 n806 3 1 2 n808-2 n809-2
0 n875 6 1 2 n876-1 n877-1
0 n874 3 1 2 n876-2 n877-2
2 n583-1 1 n583 
2 n583-2 1 n583 
2 n583-3 1 n583 
2 n762-1 1 n762 
2 n762-2 1 n762 
2 n762-3 1 n762 
2 n841-1 1 n841 
2 n841-2 1 n841 
0 n580 4 1 2 n583-1 n584-1
0 n582 5 2 1 n583-2
0 n587 6 1 2 n583-3 n584-2
0 n479 6 7 2 n615 n616
0 n440 6 7 2 n661 n662
0 n480 6 7 2 n705 n706
0 n759 4 1 2 n762-1 n763-1
0 n761 5 2 1 n762-2
0 n766 6 1 2 n762-3 n763-2
0 n799 7 2 2 n806 n807
0 n839 6 1 2 n840-1 n841-1
0 n838 3 1 2 n840-2 n841-2
0 n425 6 8 2 n874 n875
0 n433 6 7 2 n838 n839
2 n582-1 1 n582 
2 n582-2 1 n582 
2 n479-1 1 n479 
2 n479-2 1 n479 
2 n479-3 1 n479 
2 n479-4 1 n479 
2 n479-5 1 n479 
2 n479-6 1 n479 
2 n479-7 1 n479 
2 n440-1 1 n440 
2 n440-2 1 n440 
2 n440-3 1 n440 
2 n440-4 1 n440 
2 n440-5 1 n440 
2 n440-6 1 n440 
2 n440-7 1 n440 
2 n480-1 1 n480 
2 n480-2 1 n480 
2 n480-3 1 n480 
2 n480-4 1 n480 
2 n480-5 1 n480 
2 n480-6 1 n480 
2 n480-7 1 n480 
2 n761-1 1 n761 
2 n761-2 1 n761 
2 n799-1 1 n799 
2 n799-2 1 n799 
2 n425-1 1 n425 
2 n425-2 1 n425 
2 n425-3 1 n425 
2 n425-4 1 n425 
2 n425-5 1 n425 
2 n425-6 1 n425 
2 n425-7 1 n425 
2 n425-8 1 n425 
0 n474 4 1 2 n479-1 n480-1
0 n502 5 2 1 n425-5
0 n581 4 1 2 N69-3 n582-1
0 n588 6 1 2 N69-4 n582-2
0 n456 5 3 1 n440-6
0 n459 5 2 1 n480-6
0 n441 5 4 1 n479-7
0 n506 4 3 2 n440-7 n480-7
0 n760 4 1 2 N1-3 n761-1
0 n767 6 1 2 N1-4 n761-2
0 n797 6 1 2 n798-1 n799-1
0 n796 3 1 2 n798-2 n799-2
2 n433-1 1 n433 
2 n433-2 1 n433 
2 n433-3 1 n433 
2 n433-4 1 n433 
2 n433-5 1 n433 
2 n433-6 1 n433 
2 n433-7 1 n433 
0 n503 5 2 1 n433-5
0 n574 4 1 2 n580 n581
0 n586 6 1 2 n587 n588
0 n754 4 1 2 n759 n760
0 n765 6 1 2 n766 n767
0 n499 6 3 2 n796 n797
0 n505 4 3 2 n433-7 n425-8
2 n502-1 1 n502 
2 n502-2 1 n502 
2 n456-1 1 n456 
2 n456-2 1 n456 
2 n456-3 1 n456 
2 n459-1 1 n459 
2 n459-2 1 n459 
2 n441-1 1 n441 
2 n441-2 1 n441 
2 n441-3 1 n441 
2 n441-4 1 n441 
2 n506-1 1 n506 
2 n506-2 1 n506 
2 n506-3 1 n506 
0 n438 6 1 2 n441-1 n440-1
0 n494 7 1 2 n479-2 n506-1
0 n573 6 1 2 n574 n575
0 n572 6 1 2 n585 n586
0 n614 4 1 2 n456-3 n459-2
0 n613 4 1 2 n441-3 n506-2
0 n569 6 1 2 n441-4 n506-3
0 n753 6 1 2 n754 n755
0 n752 6 1 2 n764 n765
2 n503-1 1 n503 
2 n503-2 1 n503 
2 n499-1 1 n499 
2 n499-2 1 n499 
2 n499-3 1 n499 
2 n505-1 1 n505 
2 n505-2 1 n505 
2 n505-3 1 n505 
0 n501 4 1 2 n502-1 n503-1
0 n478 6 6 2 n572 n573
0 n571 4 1 2 n613 n614
0 n429 6 8 2 n752 n753
0 n437 5 6 1 n499-3
2 n478-1 1 n478 
2 n478-2 1 n478 
2 n478-3 1 n478 
2 n478-4 1 n478 
2 n478-5 1 n478 
2 n478-6 1 n478 
2 n429-1 1 n429 
2 n429-2 1 n429 
2 n429-3 1 n429 
2 n429-4 1 n429 
2 n429-5 1 n429 
2 n429-6 1 n429 
2 n429-7 1 n429 
2 n429-8 1 n429 
2 n437-1 1 n437 
2 n437-2 1 n437 
2 n437-3 1 n437 
2 n437-4 1 n437 
2 n437-5 1 n437 
2 n437-6 1 n437 
0 n520 4 1 2 n502-2 n429-5
0 n536 4 1 2 n503-2 n437-5
0 n504 5 3 1 n429-6
0 n551 4 1 2 n429-7 n499-2
0 n458 5 3 1 n478-6
0 n567 7 1 2 n437-6 n505-3
2 n504-1 1 n504 
2 n504-2 1 n504 
2 n504-3 1 n504 
2 n458-1 1 n458 
2 n458-2 1 n458 
2 n458-3 1 n458 
0 n500 4 1 2 n504-1 n505-1
0 n496 6 1 2 n504-2 n505-2
0 n535 4 1 2 n504-3 n425-6
0 n570 6 1 2 n571 n458-3
0 n498 4 1 2 n500 n501
0 n537 6 3 2 n569 n570
0 n497 6 1 2 n498 n499-1
2 n537-1 1 n537 
2 n537-2 1 n537 
2 n537-3 1 n537 
0 n477 6 2 2 n496 n497
0 n521 7 2 2 n536 n537-1
0 n553 6 1 2 n537-2 n425-7
0 n568 7 1 2 n537-3 n429-8
0 n552 4 1 2 n553 n433-6
0 n557 7 4 2 n567 n568
2 n477-1 1 n477 
2 n477-2 1 n477 
2 n521-1 1 n521 
2 n521-2 1 n521 
0 n476 6 1 2 n477-1 n478-1
0 n460 5 2 1 n477-2
0 n510 7 4 2 n520 n521-1
0 n525 7 4 2 n535 n521-2
0 n541 7 4 2 n551 n552
2 n557-1 1 n557 
2 n557-2 1 n557 
2 n557-3 1 n557 
2 n557-4 1 n557 
0 n475 4 1 2 n476 n456-2
0 n556 6 2 2 n557-1 n440-5
0 n560 6 2 2 n557-2 n479-6
0 n563 6 2 2 n557-3 n480-5
0 n566 6 2 2 n557-4 n478-5
2 n460-1 1 n460 
2 n460-2 1 n460 
2 n510-1 1 n510 
2 n510-2 1 n510 
2 n510-3 1 n510 
2 n510-4 1 n510 
2 n525-1 1 n525 
2 n525-2 1 n525 
2 n525-3 1 n525 
2 n525-4 1 n525 
2 n541-1 1 n541 
2 n541-2 1 n541 
2 n541-3 1 n541 
2 n541-4 1 n541 
0 n457 4 1 2 n460-1 n459-1
0 n464 7 4 2 n474 n475
0 n495 4 1 2 n460-2 n458-2
0 n509 6 2 2 n510-1 n440-2
0 n513 6 2 2 n510-2 n479-3
0 n516 6 2 2 n510-3 n480-2
0 n519 6 2 2 n510-4 n478-2
0 n524 6 2 2 n525-1 n440-3
0 n528 6 2 2 n525-2 n479-4
0 n531 6 2 2 n525-3 n480-3
0 n534 6 2 2 n525-4 n478-3
0 n540 6 2 2 n541-1 n440-4
0 n544 6 2 2 n541-2 n479-5
0 n547 6 2 2 n541-3 n480-4
0 n550 6 2 2 n541-4 n478-4
2 n556-1 1 n556 
2 n556-2 1 n556 
2 n560-1 1 n560 
2 n560-2 1 n560 
2 n563-1 1 n563 
2 n563-2 1 n563 
2 n566-1 1 n566 
2 n566-2 1 n566 
0 n439 6 2 2 n457 n458-1
0 n484 7 4 2 n494 n495
0 n555 6 1 2 N13-1 n556-1
0 n554 3 1 2 N13-2 n556-2
0 n559 6 1 2 N9-1 n560-1
0 n558 3 1 2 N9-2 n560-2
0 n562 6 1 2 N5-1 n563-1
0 n561 3 1 2 N5-2 n563-2
0 n565 6 1 2 N1-1 n566-1
0 n564 3 1 2 N1-2 n566-2
2 n464-1 1 n464 
2 n464-2 1 n464 
2 n464-3 1 n464 
2 n464-4 1 n464 
2 n509-1 1 n509 
2 n509-2 1 n509 
2 n513-1 1 n513 
2 n513-2 1 n513 
2 n516-1 1 n516 
2 n516-2 1 n516 
2 n519-1 1 n519 
2 n519-2 1 n519 
2 n524-1 1 n524 
2 n524-2 1 n524 
2 n528-1 1 n528 
2 n528-2 1 n528 
2 n531-1 1 n531 
2 n531-2 1 n531 
2 n534-1 1 n534 
2 n534-2 1 n534 
2 n540-1 1 n540 
2 n540-2 1 n540 
2 n544-1 1 n544 
2 n544-2 1 n544 
2 n547-1 1 n547 
2 n547-2 1 n547 
2 n550-1 1 n550 
2 n550-2 1 n550 
0 n463 6 2 2 n464-1 n425-3
0 n467 6 2 2 n464-2 n429-3
0 n470 6 2 2 n464-3 n433-3
0 n473 6 2 2 n464-4 n437-3
0 n508 6 1 2 N61-1 n509-1
0 n507 3 1 2 N61-2 n509-2
0 n512 6 1 2 N57-1 n513-1
0 n511 3 1 2 N57-2 n513-2
0 n515 6 1 2 N53-1 n516-1
0 n514 3 1 2 N53-2 n516-2
0 n518 6 1 2 N49-1 n519-1
0 n517 3 1 2 N49-2 n519-2
0 n523 6 1 2 N45-1 n524-1
0 n522 3 1 2 N45-2 n524-2
0 n527 6 1 2 N41-1 n528-1
0 n526 3 1 2 N41-2 n528-2
0 n530 6 1 2 N37-1 n531-1
0 n529 3 1 2 N37-2 n531-2
0 n533 6 1 2 N33-1 n534-1
0 n532 3 1 2 N33-2 n534-2
0 n539 6 1 2 N29-1 n540-1
0 n538 3 1 2 N29-2 n540-2
0 n543 6 1 2 N25-1 n544-1
0 n542 3 1 2 N25-2 n544-2
0 n546 6 1 2 N21-1 n547-1
0 n545 3 1 2 N21-2 n547-2
0 n549 6 1 2 N17-1 n550-1
0 n548 3 1 2 N17-2 n550-2
3 N727 6 0 2 n554 n555
3 N726 6 0 2 n558 n559
3 N725 6 0 2 n561 n562
3 N724 6 0 2 n564 n565
2 n439-1 1 n439 
2 n439-2 1 n439 
2 n484-1 1 n484 
2 n484-2 1 n484 
2 n484-3 1 n484 
2 n484-4 1 n484 
0 n424 4 4 2 n438 n439-1
0 n455 4 1 2 n439-2 n441-2
0 n483 6 2 2 n484-1 n425-4
0 n487 6 2 2 n484-2 n429-4
0 n490 6 2 2 n484-3 n433-4
0 n493 6 2 2 n484-4 n437-4
3 N739 6 0 2 n507 n508
3 N738 6 0 2 n511 n512
3 N737 6 0 2 n514 n515
3 N736 6 0 2 n517 n518
3 N735 6 0 2 n522 n523
3 N734 6 0 2 n526 n527
3 N733 6 0 2 n529 n530
3 N732 6 0 2 n532 n533
3 N731 6 0 2 n538 n539
3 N730 6 0 2 n542 n543
3 N729 6 0 2 n545 n546
3 N728 6 0 2 n548 n549
2 n463-1 1 n463 
2 n463-2 1 n463 
2 n467-1 1 n467 
2 n467-2 1 n467 
2 n470-1 1 n470 
2 n470-2 1 n470 
2 n473-1 1 n473 
2 n473-2 1 n473 
0 n445 7 4 2 n455 n456-1
0 n462 6 1 2 N93-1 n463-1
0 n461 3 1 2 N93-2 n463-2
0 n466 6 1 2 N89-1 n467-1
0 n465 3 1 2 N89-2 n467-2
0 n469 6 1 2 N85-1 n470-1
0 n468 3 1 2 N85-2 n470-2
0 n472 6 1 2 N81-1 n473-1
0 n471 3 1 2 N81-2 n473-2
2 n424-1 1 n424 
2 n424-2 1 n424 
2 n424-3 1 n424 
2 n424-4 1 n424 
2 n483-1 1 n483 
2 n483-2 1 n483 
2 n487-1 1 n487 
2 n487-2 1 n487 
2 n490-1 1 n490 
2 n490-2 1 n490 
2 n493-1 1 n493 
2 n493-2 1 n493 
0 n423 6 2 2 n424-1 n425-1
0 n428 6 2 2 n424-2 n429-1
0 n432 6 2 2 n424-3 n433-1
0 n436 6 2 2 n424-4 n437-1
3 N747 6 0 2 n461 n462
3 N746 6 0 2 n465 n466
3 N745 6 0 2 n468 n469
3 N744 6 0 2 n471 n472
0 n482 6 1 2 N77-1 n483-1
0 n481 3 1 2 N77-2 n483-2
0 n486 6 1 2 N73-1 n487-1
0 n485 3 1 2 N73-2 n487-2
0 n489 6 1 2 N69-1 n490-1
0 n488 3 1 2 N69-2 n490-2
0 n492 6 1 2 N65-1 n493-1
0 n491 3 1 2 N65-2 n493-2
2 n445-1 1 n445 
2 n445-2 1 n445 
2 n445-3 1 n445 
2 n445-4 1 n445 
0 n444 6 2 2 n445-1 n425-2
0 n448 6 2 2 n445-2 n429-2
0 n451 6 2 2 n445-3 n433-2
0 n454 6 2 2 n445-4 n437-2
3 N743 6 0 2 n481 n482
3 N742 6 0 2 n485 n486
3 N741 6 0 2 n488 n489
3 N740 6 0 2 n491 n492
2 n423-1 1 n423 
2 n423-2 1 n423 
2 n428-1 1 n428 
2 n428-2 1 n428 
2 n432-1 1 n432 
2 n432-2 1 n432 
2 n436-1 1 n436 
2 n436-2 1 n436 
0 n422 6 1 2 N125-1 n423-1
0 n421 3 1 2 N125-2 n423-2
0 n427 6 1 2 N121-1 n428-1
0 n426 3 1 2 N121-2 n428-2
0 n431 6 1 2 N117-1 n432-1
0 n430 3 1 2 N117-2 n432-2
0 n435 6 1 2 N113-1 n436-1
0 n434 3 1 2 N113-2 n436-2
2 n444-1 1 n444 
2 n444-2 1 n444 
2 n448-1 1 n448 
2 n448-2 1 n448 
2 n451-1 1 n451 
2 n451-2 1 n451 
2 n454-1 1 n454 
2 n454-2 1 n454 
3 N755 6 0 2 n421 n422
3 N754 6 0 2 n426 n427
3 N753 6 0 2 n430 n431
3 N752 6 0 2 n434 n435
0 n443 6 1 2 N109-1 n444-1
0 n442 3 1 2 N109-2 n444-2
0 n447 6 1 2 N105-1 n448-1
0 n446 3 1 2 N105-2 n448-2
0 n450 6 1 2 N101-1 n451-1
0 n449 3 1 2 N101-2 n451-2
0 n453 6 1 2 N97-1 n454-1
0 n452 3 1 2 N97-2 n454-2
3 N751 6 0 2 n442 n443
3 N750 6 0 2 n446 n447
3 N749 6 0 2 n449 n450
3 N748 6 0 2 n452 n453
