1	1	0	16	0	
1	18	0	16	0	
1	35	0	16	0	
1	52	0	16	0	
1	69	0	16	0	
1	86	0	16	0	
1	103	0	16	0	
1	120	0	16	0	
1	137	0	16	0	
1	154	0	16	0	
1	171	0	16	0	
1	188	0	16	0	
1	205	0	16	0	
1	222	0	16	0	
1	239	0	16	0	
1	256	0	16	0	
1	273	0	16	0	
1	290	0	16	0	
1	307	0	16	0	
1	324	0	16	0	
1	341	0	16	0	
1	358	0	16	0	
1	375	0	16	0	
1	392	0	16	0	
1	409	0	16	0	
1	426	0	16	0	
1	443	0	16	0	
1	460	0	16	0	
1	477	0	16	0	
1	494	0	16	0	
1	511	0	16	0	
1	528	0	16	0	
3	545	7	0	2	6289	6545	
0	546	7	2	2	6290	6561	
0	549	7	2	2	6291	6577	
0	552	7	2	2	6292	6593	
0	555	7	2	2	6293	6609	
0	558	7	2	2	6294	6625	
0	561	7	2	2	6295	6641	
0	564	7	2	2	6296	6657	
0	567	7	2	2	6297	6673	
0	570	7	2	2	6298	6689	
0	573	7	2	2	6299	6705	
0	576	7	2	2	6300	6721	
0	579	7	2	2	6301	6737	
0	582	7	2	2	6302	6753	
0	585	7	2	2	6303	6769	
0	588	7	2	2	6304	6785	
0	591	7	2	2	6305	6546	
0	594	7	2	2	6306	6562	
0	597	7	2	2	6307	6578	
0	600	7	2	2	6308	6594	
0	603	7	2	2	6309	6610	
0	606	7	2	2	6310	6626	
0	609	7	2	2	6311	6642	
0	612	7	2	2	6312	6658	
0	615	7	2	2	6313	6674	
0	618	7	2	2	6314	6690	
0	621	7	2	2	6315	6706	
0	624	7	2	2	6316	6722	
0	627	7	2	2	6317	6738	
0	630	7	2	2	6318	6754	
0	633	7	2	2	6319	6770	
0	636	7	2	2	6320	6786	
0	639	7	2	2	6321	6547	
0	642	7	2	2	6322	6563	
0	645	7	2	2	6323	6579	
0	648	7	2	2	6324	6595	
0	651	7	2	2	6325	6611	
0	654	7	2	2	6326	6627	
0	657	7	2	2	6327	6643	
0	660	7	2	2	6328	6659	
0	663	7	2	2	6329	6675	
0	666	7	2	2	6330	6691	
0	669	7	2	2	6331	6707	
0	672	7	2	2	6332	6723	
0	675	7	2	2	6333	6739	
0	678	7	2	2	6334	6755	
0	681	7	2	2	6335	6771	
0	684	7	2	2	6336	6787	
0	687	7	2	2	6337	6548	
0	690	7	2	2	6338	6564	
0	693	7	2	2	6339	6580	
0	696	7	2	2	6340	6596	
0	699	7	2	2	6341	6612	
0	702	7	2	2	6342	6628	
0	705	7	2	2	6343	6644	
0	708	7	2	2	6344	6660	
0	711	7	2	2	6345	6676	
0	714	7	2	2	6346	6692	
0	717	7	2	2	6347	6708	
0	720	7	2	2	6348	6724	
0	723	7	2	2	6349	6740	
0	726	7	2	2	6350	6756	
0	729	7	2	2	6351	6772	
0	732	7	2	2	6352	6788	
0	735	7	2	2	6353	6549	
0	738	7	2	2	6354	6565	
0	741	7	2	2	6355	6581	
0	744	7	2	2	6356	6597	
0	747	7	2	2	6357	6613	
0	750	7	2	2	6358	6629	
0	753	7	2	2	6359	6645	
0	756	7	2	2	6360	6661	
0	759	7	2	2	6361	6677	
0	762	7	2	2	6362	6693	
0	765	7	2	2	6363	6709	
0	768	7	2	2	6364	6725	
0	771	7	2	2	6365	6741	
0	774	7	2	2	6366	6757	
0	777	7	2	2	6367	6773	
0	780	7	2	2	6368	6789	
0	783	7	2	2	6369	6550	
0	786	7	2	2	6370	6566	
0	789	7	2	2	6371	6582	
0	792	7	2	2	6372	6598	
0	795	7	2	2	6373	6614	
0	798	7	2	2	6374	6630	
0	801	7	2	2	6375	6646	
0	804	7	2	2	6376	6662	
0	807	7	2	2	6377	6678	
0	810	7	2	2	6378	6694	
0	813	7	2	2	6379	6710	
0	816	7	2	2	6380	6726	
0	819	7	2	2	6381	6742	
0	822	7	2	2	6382	6758	
0	825	7	2	2	6383	6774	
0	828	7	2	2	6384	6790	
0	831	7	2	2	6385	6551	
0	834	7	2	2	6386	6567	
0	837	7	2	2	6387	6583	
0	840	7	2	2	6388	6599	
0	843	7	2	2	6389	6615	
0	846	7	2	2	6390	6631	
0	849	7	2	2	6391	6647	
0	852	7	2	2	6392	6663	
0	855	7	2	2	6393	6679	
0	858	7	2	2	6394	6695	
0	861	7	2	2	6395	6711	
0	864	7	2	2	6396	6727	
0	867	7	2	2	6397	6743	
0	870	7	2	2	6398	6759	
0	873	7	2	2	6399	6775	
0	876	7	2	2	6400	6791	
0	879	7	2	2	6401	6552	
0	882	7	2	2	6402	6568	
0	885	7	2	2	6403	6584	
0	888	7	2	2	6404	6600	
0	891	7	2	2	6405	6616	
0	894	7	2	2	6406	6632	
0	897	7	2	2	6407	6648	
0	900	7	2	2	6408	6664	
0	903	7	2	2	6409	6680	
0	906	7	2	2	6410	6696	
0	909	7	2	2	6411	6712	
0	912	7	2	2	6412	6728	
0	915	7	2	2	6413	6744	
0	918	7	2	2	6414	6760	
0	921	7	2	2	6415	6776	
0	924	7	2	2	6416	6792	
0	927	7	2	2	6417	6553	
0	930	7	2	2	6418	6569	
0	933	7	2	2	6419	6585	
0	936	7	2	2	6420	6601	
0	939	7	2	2	6421	6617	
0	942	7	2	2	6422	6633	
0	945	7	2	2	6423	6649	
0	948	7	2	2	6424	6665	
0	951	7	2	2	6425	6681	
0	954	7	2	2	6426	6697	
0	957	7	2	2	6427	6713	
0	960	7	2	2	6428	6729	
0	963	7	2	2	6429	6745	
0	966	7	2	2	6430	6761	
0	969	7	2	2	6431	6777	
0	972	7	2	2	6432	6793	
0	975	7	2	2	6433	6554	
0	978	7	2	2	6434	6570	
0	981	7	2	2	6435	6586	
0	984	7	2	2	6436	6602	
0	987	7	2	2	6437	6618	
0	990	7	2	2	6438	6634	
0	993	7	2	2	6439	6650	
0	996	7	2	2	6440	6666	
0	999	7	2	2	6441	6682	
0	1002	7	2	2	6442	6698	
0	1005	7	2	2	6443	6714	
0	1008	7	2	2	6444	6730	
0	1011	7	2	2	6445	6746	
0	1014	7	2	2	6446	6762	
0	1017	7	2	2	6447	6778	
0	1020	7	2	2	6448	6794	
0	1023	7	2	2	6449	6555	
0	1026	7	2	2	6450	6571	
0	1029	7	2	2	6451	6587	
0	1032	7	2	2	6452	6603	
0	1035	7	2	2	6453	6619	
0	1038	7	2	2	6454	6635	
0	1041	7	2	2	6455	6651	
0	1044	7	2	2	6456	6667	
0	1047	7	2	2	6457	6683	
0	1050	7	2	2	6458	6699	
0	1053	7	2	2	6459	6715	
0	1056	7	2	2	6460	6731	
0	1059	7	2	2	6461	6747	
0	1062	7	2	2	6462	6763	
0	1065	7	2	2	6463	6779	
0	1068	7	2	2	6464	6795	
0	1071	7	2	2	6465	6556	
0	1074	7	2	2	6466	6572	
0	1077	7	2	2	6467	6588	
0	1080	7	2	2	6468	6604	
0	1083	7	2	2	6469	6620	
0	1086	7	2	2	6470	6636	
0	1089	7	2	2	6471	6652	
0	1092	7	2	2	6472	6668	
0	1095	7	2	2	6473	6684	
0	1098	7	2	2	6474	6700	
0	1101	7	2	2	6475	6716	
0	1104	7	2	2	6476	6732	
0	1107	7	2	2	6477	6748	
0	1110	7	2	2	6478	6764	
0	1113	7	2	2	6479	6780	
0	1116	7	2	2	6480	6796	
0	1119	7	2	2	6481	6557	
0	1122	7	2	2	6482	6573	
0	1125	7	2	2	6483	6589	
0	1128	7	2	2	6484	6605	
0	1131	7	2	2	6485	6621	
0	1134	7	2	2	6486	6637	
0	1137	7	2	2	6487	6653	
0	1140	7	2	2	6488	6669	
0	1143	7	2	2	6489	6685	
0	1146	7	2	2	6490	6701	
0	1149	7	2	2	6491	6717	
0	1152	7	2	2	6492	6733	
0	1155	7	2	2	6493	6749	
0	1158	7	2	2	6494	6765	
0	1161	7	2	2	6495	6781	
0	1164	7	2	2	6496	6797	
0	1167	7	2	2	6497	6558	
0	1170	7	2	2	6498	6574	
0	1173	7	2	2	6499	6590	
0	1176	7	2	2	6500	6606	
0	1179	7	2	2	6501	6622	
0	1182	7	2	2	6502	6638	
0	1185	7	2	2	6503	6654	
0	1188	7	2	2	6504	6670	
0	1191	7	2	2	6505	6686	
0	1194	7	2	2	6506	6702	
0	1197	7	2	2	6507	6718	
0	1200	7	2	2	6508	6734	
0	1203	7	2	2	6509	6750	
0	1206	7	2	2	6510	6766	
0	1209	7	2	2	6511	6782	
0	1212	7	2	2	6512	6798	
0	1215	7	2	2	6513	6559	
0	1218	7	2	2	6514	6575	
0	1221	7	2	2	6515	6591	
0	1224	7	2	2	6516	6607	
0	1227	7	2	2	6517	6623	
0	1230	7	2	2	6518	6639	
0	1233	7	2	2	6519	6655	
0	1236	7	2	2	6520	6671	
0	1239	7	2	2	6521	6687	
0	1242	7	2	2	6522	6703	
0	1245	7	2	2	6523	6719	
0	1248	7	2	2	6524	6735	
0	1251	7	2	2	6525	6751	
0	1254	7	2	2	6526	6767	
0	1257	7	2	2	6527	6783	
0	1260	7	2	2	6528	6799	
0	1263	7	2	2	6529	6560	
0	1266	7	2	2	6530	6576	
0	1269	7	2	2	6531	6592	
0	1272	7	2	2	6532	6608	
0	1275	7	2	2	6533	6624	
0	1278	7	2	2	6534	6640	
0	1281	7	2	2	6535	6656	
0	1284	7	2	2	6536	6672	
0	1287	7	2	2	6537	6688	
0	1290	7	2	2	6538	6704	
0	1293	7	2	2	6539	6720	
0	1296	7	2	2	6540	6736	
0	1299	7	2	2	6541	6752	
0	1302	7	2	2	6542	6768	
0	1305	7	2	2	6543	6784	
0	1308	7	2	2	6544	6800	
0	1311	5	3	1	6831	
0	1315	5	3	1	6863	
0	1319	5	3	1	6895	
0	1323	5	3	1	6927	
0	1327	5	3	1	6959	
0	1331	5	3	1	6991	
0	1335	5	3	1	7023	
0	1339	5	3	1	7055	
0	1343	5	3	1	7087	
0	1347	5	3	1	7119	
0	1351	5	3	1	7151	
0	1355	5	3	1	7183	
0	1359	5	3	1	7215	
0	1363	5	3	1	7247	
0	1367	5	3	1	7279	
0	1371	4	1	2	6832	7311	
0	1372	5	1	1	7312	
0	1373	4	1	2	6864	7314	
0	1374	5	1	1	7315	
0	1375	4	1	2	6896	7317	
0	1376	5	1	1	7318	
0	1377	4	1	2	6928	7320	
0	1378	5	1	1	7321	
0	1379	4	1	2	6960	7323	
0	1380	5	1	1	7324	
0	1381	4	1	2	6992	7326	
0	1382	5	1	1	7327	
0	1383	4	1	2	7024	7329	
0	1384	5	1	1	7330	
0	1385	4	1	2	7056	7332	
0	1386	5	1	1	7333	
0	1387	4	1	2	7088	7335	
0	1388	5	1	1	7336	
0	1389	4	1	2	7120	7338	
0	1390	5	1	1	7339	
0	1391	4	1	2	7152	7341	
0	1392	5	1	1	7342	
0	1393	4	1	2	7184	7344	
0	1394	5	1	1	7345	
0	1395	4	1	2	7216	7347	
0	1396	5	1	1	7348	
0	1397	4	1	2	7248	7350	
0	1398	5	1	1	7351	
0	1399	4	1	2	7280	7353	
0	1400	5	1	1	7354	
0	1401	4	2	2	1371	1372	
0	1404	4	2	2	1373	1374	
0	1407	4	2	2	1375	1376	
0	1410	4	2	2	1377	1378	
0	1413	4	2	2	1379	1380	
0	1416	4	2	2	1381	1382	
0	1419	4	2	2	1383	1384	
0	1422	4	2	2	1385	1386	
0	1425	4	2	2	1387	1388	
0	1428	4	2	2	1389	1390	
0	1431	4	2	2	1391	1392	
0	1434	4	2	2	1393	1394	
0	1437	4	2	2	1395	1396	
0	1440	4	2	2	1397	1398	
0	1443	4	2	2	1399	1400	
0	1446	4	3	2	7356	6801	
0	1450	4	3	2	7358	6833	
0	1454	4	3	2	7360	6865	
0	1458	4	3	2	7362	6897	
0	1462	4	3	2	7364	6929	
0	1466	4	3	2	7366	6961	
0	1470	4	3	2	7368	6993	
0	1474	4	3	2	7370	7025	
0	1478	4	3	2	7372	7057	
0	1482	4	3	2	7374	7089	
0	1486	4	3	2	7376	7121	
0	1490	4	3	2	7378	7153	
0	1494	4	3	2	7380	7185	
0	1498	4	3	2	7382	7217	
0	1502	4	3	2	7384	7249	
0	1506	4	1	2	7357	7386	
0	1507	4	1	2	7387	6802	
0	1508	4	2	2	7313	7388	
0	1511	4	1	2	7359	7389	
0	1512	4	1	2	7390	6834	
0	1513	4	2	2	7316	7391	
0	1516	4	1	2	7361	7392	
0	1517	4	1	2	7393	6866	
0	1518	4	2	2	7319	7394	
0	1521	4	1	2	7363	7395	
0	1522	4	1	2	7396	6898	
0	1523	4	2	2	7322	7397	
0	1526	4	1	2	7365	7398	
0	1527	4	1	2	7399	6930	
0	1528	4	2	2	7325	7400	
0	1531	4	1	2	7367	7401	
0	1532	4	1	2	7402	6962	
0	1533	4	2	2	7328	7403	
0	1536	4	1	2	7369	7404	
0	1537	4	1	2	7405	6994	
0	1538	4	2	2	7331	7406	
0	1541	4	1	2	7371	7407	
0	1542	4	1	2	7408	7026	
0	1543	4	2	2	7334	7409	
0	1546	4	1	2	7373	7410	
0	1547	4	1	2	7411	7058	
0	1548	4	2	2	7337	7412	
0	1551	4	1	2	7375	7413	
0	1552	4	1	2	7414	7090	
0	1553	4	2	2	7340	7415	
0	1556	4	1	2	7377	7416	
0	1557	4	1	2	7417	7122	
0	1558	4	2	2	7343	7418	
0	1561	4	1	2	7379	7419	
0	1562	4	1	2	7420	7154	
0	1563	4	2	2	7346	7421	
0	1566	4	1	2	7381	7422	
0	1567	4	1	2	7423	7186	
0	1568	4	2	2	7349	7424	
0	1571	4	1	2	7383	7425	
0	1572	4	1	2	7426	7218	
0	1573	4	2	2	7352	7427	
0	1576	4	1	2	7385	7428	
0	1577	4	1	2	7429	7250	
0	1578	4	2	2	7355	7430	
3	1581	4	0	2	1506	1507	
0	1582	4	2	2	1511	1512	
0	1585	4	2	2	1516	1517	
0	1588	4	2	2	1521	1522	
0	1591	4	2	2	1526	1527	
0	1594	4	2	2	1531	1532	
0	1597	4	2	2	1536	1537	
0	1600	4	2	2	1541	1542	
0	1603	4	2	2	1546	1547	
0	1606	4	2	2	1551	1552	
0	1609	4	2	2	1556	1557	
0	1612	4	2	2	1561	1562	
0	1615	4	2	2	1566	1567	
0	1618	4	2	2	1571	1572	
0	1621	4	2	2	1576	1577	
0	1624	4	3	2	7281	7459	
0	1628	4	3	2	7461	7431	
0	1632	4	3	2	7463	7433	
0	1636	4	3	2	7465	7435	
0	1640	4	3	2	7467	7437	
0	1644	4	3	2	7469	7439	
0	1648	4	3	2	7471	7441	
0	1652	4	3	2	7473	7443	
0	1656	4	3	2	7475	7445	
0	1660	4	3	2	7477	7447	
0	1664	4	3	2	7479	7449	
0	1668	4	3	2	7481	7451	
0	1672	4	3	2	7483	7453	
0	1676	4	3	2	7485	7455	
0	1680	4	3	2	7487	7457	
0	1684	4	1	2	7282	7489	
0	1685	4	1	2	7490	7460	
0	1686	4	1	2	7462	7492	
0	1687	4	1	2	7493	7432	
0	1688	4	1	2	7464	7495	
0	1689	4	1	2	7496	7434	
0	1690	4	1	2	7466	7498	
0	1691	4	1	2	7499	7436	
0	1692	4	1	2	7468	7501	
0	1693	4	1	2	7502	7438	
0	1694	4	1	2	7470	7504	
0	1695	4	1	2	7505	7440	
0	1696	4	1	2	7472	7507	
0	1697	4	1	2	7508	7442	
0	1698	4	1	2	7474	7510	
0	1699	4	1	2	7511	7444	
0	1700	4	1	2	7476	7513	
0	1701	4	1	2	7514	7446	
0	1702	4	1	2	7478	7516	
0	1703	4	1	2	7517	7448	
0	1704	4	1	2	7480	7519	
0	1705	4	1	2	7520	7450	
0	1706	4	1	2	7482	7522	
0	1707	4	1	2	7523	7452	
0	1708	4	1	2	7484	7525	
0	1709	4	1	2	7526	7454	
0	1710	4	1	2	7486	7528	
0	1711	4	1	2	7529	7456	
0	1712	4	1	2	7488	7531	
0	1713	4	1	2	7532	7458	
0	1714	4	2	2	1684	1685	
0	1717	4	2	2	1686	1687	
0	1720	4	2	2	1688	1689	
0	1723	4	2	2	1690	1691	
0	1726	4	2	2	1692	1693	
0	1729	4	2	2	1694	1695	
0	1732	4	2	2	1696	1697	
0	1735	4	2	2	1698	1699	
0	1738	4	2	2	1700	1701	
0	1741	4	2	2	1702	1703	
0	1744	4	2	2	1704	1705	
0	1747	4	2	2	1706	1707	
0	1750	4	2	2	1708	1709	
0	1753	4	2	2	1710	1711	
0	1756	4	2	2	1712	1713	
0	1759	4	3	2	7534	7251	
0	1763	4	3	2	7536	6803	
0	1767	4	3	2	7538	6835	
0	1771	4	3	2	7540	6867	
0	1775	4	3	2	7542	6899	
0	1779	4	3	2	7544	6931	
0	1783	4	3	2	7546	6963	
0	1787	4	3	2	7548	6995	
0	1791	4	3	2	7550	7027	
0	1795	4	3	2	7552	7059	
0	1799	4	3	2	7554	7091	
0	1803	4	3	2	7556	7123	
0	1807	4	3	2	7558	7155	
0	1811	4	3	2	7560	7187	
0	1815	4	3	2	7562	7219	
0	1819	4	1	2	7535	7564	
0	1820	4	1	2	7565	7252	
0	1821	4	2	2	7491	7566	
0	1824	4	1	2	7537	7567	
0	1825	4	1	2	7568	6804	
0	1826	4	2	2	7494	7569	
0	1829	4	1	2	7539	7570	
0	1830	4	1	2	7571	6836	
0	1831	4	2	2	7497	7572	
0	1834	4	1	2	7541	7573	
0	1835	4	1	2	7574	6868	
0	1836	4	2	2	7500	7575	
0	1839	4	1	2	7543	7576	
0	1840	4	1	2	7577	6900	
0	1841	4	2	2	7503	7578	
0	1844	4	1	2	7545	7579	
0	1845	4	1	2	7580	6932	
0	1846	4	2	2	7506	7581	
0	1849	4	1	2	7547	7582	
0	1850	4	1	2	7583	6964	
0	1851	4	2	2	7509	7584	
0	1854	4	1	2	7549	7585	
0	1855	4	1	2	7586	6996	
0	1856	4	2	2	7512	7587	
0	1859	4	1	2	7551	7588	
0	1860	4	1	2	7589	7028	
0	1861	4	2	2	7515	7590	
0	1864	4	1	2	7553	7591	
0	1865	4	1	2	7592	7060	
0	1866	4	2	2	7518	7593	
0	1869	4	1	2	7555	7594	
0	1870	4	1	2	7595	7092	
0	1871	4	2	2	7521	7596	
0	1874	4	1	2	7557	7597	
0	1875	4	1	2	7598	7124	
0	1876	4	2	2	7524	7599	
0	1879	4	1	2	7559	7600	
0	1880	4	1	2	7601	7156	
0	1881	4	2	2	7527	7602	
0	1884	4	1	2	7561	7603	
0	1885	4	1	2	7604	7188	
0	1886	4	2	2	7530	7605	
0	1889	4	1	2	7563	7606	
0	1890	4	1	2	7607	7220	
0	1891	4	2	2	7533	7608	
0	1894	4	2	2	1819	1820	
0	1897	4	3	2	7283	7609	
3	1901	4	0	2	1824	1825	
0	1902	4	2	2	1829	1830	
0	1905	4	2	2	1834	1835	
0	1908	4	2	2	1839	1840	
0	1911	4	2	2	1844	1845	
0	1914	4	2	2	1849	1850	
0	1917	4	2	2	1854	1855	
0	1920	4	2	2	1859	1860	
0	1923	4	2	2	1864	1865	
0	1926	4	2	2	1869	1870	
0	1929	4	2	2	1874	1875	
0	1932	4	2	2	1879	1880	
0	1935	4	2	2	1884	1885	
0	1938	4	2	2	1889	1890	
0	1941	4	3	2	7639	7637	
0	1945	4	1	2	7284	7641	
0	1946	4	1	2	7642	7610	
0	1947	4	3	2	7644	7611	
0	1951	4	3	2	7646	7613	
0	1955	4	3	2	7648	7615	
0	1959	4	3	2	7650	7617	
0	1963	4	3	2	7652	7619	
0	1967	4	3	2	7654	7621	
0	1971	4	3	2	7656	7623	
0	1975	4	3	2	7658	7625	
0	1979	4	3	2	7660	7627	
0	1983	4	3	2	7662	7629	
0	1987	4	3	2	7664	7631	
0	1991	4	3	2	7666	7633	
0	1995	4	3	2	7668	7635	
0	1999	4	1	2	7640	7670	
0	2000	4	1	2	7671	7638	
0	2001	4	2	2	1945	1946	
0	2004	4	1	2	7645	7673	
0	2005	4	1	2	7674	7612	
0	2006	4	1	2	7647	7676	
0	2007	4	1	2	7677	7614	
0	2008	4	1	2	7649	7679	
0	2009	4	1	2	7680	7616	
0	2010	4	1	2	7651	7682	
0	2011	4	1	2	7683	7618	
0	2012	4	1	2	7653	7685	
0	2013	4	1	2	7686	7620	
0	2014	4	1	2	7655	7688	
0	2015	4	1	2	7689	7622	
0	2016	4	1	2	7657	7691	
0	2017	4	1	2	7692	7624	
0	2018	4	1	2	7659	7694	
0	2019	4	1	2	7695	7626	
0	2020	4	1	2	7661	7697	
0	2021	4	1	2	7698	7628	
0	2022	4	1	2	7663	7700	
0	2023	4	1	2	7701	7630	
0	2024	4	1	2	7665	7703	
0	2025	4	1	2	7704	7632	
0	2026	4	1	2	7667	7706	
0	2027	4	1	2	7707	7634	
0	2028	4	1	2	7669	7709	
0	2029	4	1	2	7710	7636	
0	2030	4	2	2	1999	2000	
0	2033	4	3	2	7712	7253	
0	2037	4	2	2	2004	2005	
0	2040	4	2	2	2006	2007	
0	2043	4	2	2	2008	2009	
0	2046	4	2	2	2010	2011	
0	2049	4	2	2	2012	2013	
0	2052	4	2	2	2014	2015	
0	2055	4	2	2	2016	2017	
0	2058	4	2	2	2018	2019	
0	2061	4	2	2	2020	2021	
0	2064	4	2	2	2022	2023	
0	2067	4	2	2	2024	2025	
0	2070	4	2	2	2026	2027	
0	2073	4	2	2	2028	2029	
0	2076	4	3	2	7714	7221	
0	2080	4	1	2	7713	7716	
0	2081	4	1	2	7717	7254	
0	2082	4	2	2	7643	7718	
0	2085	4	3	2	7719	6805	
0	2089	4	3	2	7721	6837	
0	2093	4	3	2	7723	6869	
0	2097	4	3	2	7725	6901	
0	2101	4	3	2	7727	6933	
0	2105	4	3	2	7729	6965	
0	2109	4	3	2	7731	6997	
0	2113	4	3	2	7733	7029	
0	2117	4	3	2	7735	7061	
0	2121	4	3	2	7737	7093	
0	2125	4	3	2	7739	7125	
0	2129	4	3	2	7741	7157	
0	2133	4	3	2	7743	7189	
0	2137	4	1	2	7715	7745	
0	2138	4	1	2	7746	7222	
0	2139	4	2	2	7672	7747	
0	2142	4	2	2	2080	2081	
0	2145	4	3	2	7285	7748	
0	2149	4	1	2	7720	7750	
0	2150	4	1	2	7751	6806	
0	2151	4	2	2	7675	7752	
0	2154	4	1	2	7722	7753	
0	2155	4	1	2	7754	6838	
0	2156	4	2	2	7678	7755	
0	2159	4	1	2	7724	7756	
0	2160	4	1	2	7757	6870	
0	2161	4	2	2	7681	7758	
0	2164	4	1	2	7726	7759	
0	2165	4	1	2	7760	6902	
0	2166	4	2	2	7684	7761	
0	2169	4	1	2	7728	7762	
0	2170	4	1	2	7763	6934	
0	2171	4	2	2	7687	7764	
0	2174	4	1	2	7730	7765	
0	2175	4	1	2	7766	6966	
0	2176	4	2	2	7690	7767	
0	2179	4	1	2	7732	7768	
0	2180	4	1	2	7769	6998	
0	2181	4	2	2	7693	7770	
0	2184	4	1	2	7734	7771	
0	2185	4	1	2	7772	7030	
0	2186	4	2	2	7696	7773	
0	2189	4	1	2	7736	7774	
0	2190	4	1	2	7775	7062	
0	2191	4	2	2	7699	7776	
0	2194	4	1	2	7738	7777	
0	2195	4	1	2	7778	7094	
0	2196	4	2	2	7702	7779	
0	2199	4	1	2	7740	7780	
0	2200	4	1	2	7781	7126	
0	2201	4	2	2	7705	7782	
0	2204	4	1	2	7742	7783	
0	2205	4	1	2	7784	7158	
0	2206	4	2	2	7708	7785	
0	2209	4	1	2	7744	7786	
0	2210	4	1	2	7787	7190	
0	2211	4	2	2	7711	7788	
0	2214	4	2	2	2137	2138	
0	2217	4	3	2	7791	7789	
0	2221	4	1	2	7286	7793	
0	2222	4	1	2	7794	7749	
3	2223	4	0	2	2149	2150	
0	2224	4	2	2	2154	2155	
0	2227	4	2	2	2159	2160	
0	2230	4	2	2	2164	2165	
0	2233	4	2	2	2169	2170	
0	2236	4	2	2	2174	2175	
0	2239	4	2	2	2179	2180	
0	2242	4	2	2	2184	2185	
0	2245	4	2	2	2189	2190	
0	2248	4	2	2	2194	2195	
0	2251	4	2	2	2199	2200	
0	2254	4	2	2	2204	2205	
0	2257	4	2	2	2209	2210	
0	2260	4	3	2	7822	7820	
0	2264	4	1	2	7792	7824	
0	2265	4	1	2	7825	7790	
0	2266	4	2	2	2221	2222	
0	2269	4	3	2	7827	7796	
0	2273	4	3	2	7829	7798	
0	2277	4	3	2	7831	7800	
0	2281	4	3	2	7833	7802	
0	2285	4	3	2	7835	7804	
0	2289	4	3	2	7837	7806	
0	2293	4	3	2	7839	7808	
0	2297	4	3	2	7841	7810	
0	2301	4	3	2	7843	7812	
0	2305	4	3	2	7845	7814	
0	2309	4	3	2	7847	7816	
0	2313	4	3	2	7849	7818	
0	2317	4	1	2	7823	7851	
0	2318	4	1	2	7852	7821	
0	2319	4	2	2	2264	2265	
0	2322	4	3	2	7854	7255	
0	2326	4	1	2	7828	7856	
0	2327	4	1	2	7857	7797	
0	2328	4	1	2	7830	7859	
0	2329	4	1	2	7860	7799	
0	2330	4	1	2	7832	7862	
0	2331	4	1	2	7863	7801	
0	2332	4	1	2	7834	7865	
0	2333	4	1	2	7866	7803	
0	2334	4	1	2	7836	7868	
0	2335	4	1	2	7869	7805	
0	2336	4	1	2	7838	7871	
0	2337	4	1	2	7872	7807	
0	2338	4	1	2	7840	7874	
0	2339	4	1	2	7875	7809	
0	2340	4	1	2	7842	7877	
0	2341	4	1	2	7878	7811	
0	2342	4	1	2	7844	7880	
0	2343	4	1	2	7881	7813	
0	2344	4	1	2	7846	7883	
0	2345	4	1	2	7884	7815	
0	2346	4	1	2	7848	7886	
0	2347	4	1	2	7887	7817	
0	2348	4	1	2	7850	7889	
0	2349	4	1	2	7890	7819	
0	2350	4	2	2	2317	2318	
0	2353	4	3	2	7892	7223	
0	2357	4	1	2	7855	7894	
0	2358	4	1	2	7895	7256	
0	2359	4	2	2	7795	7896	
0	2362	4	2	2	2326	2327	
0	2365	4	2	2	2328	2329	
0	2368	4	2	2	2330	2331	
0	2371	4	2	2	2332	2333	
0	2374	4	2	2	2334	2335	
0	2377	4	2	2	2336	2337	
0	2380	4	2	2	2338	2339	
0	2383	4	2	2	2340	2341	
0	2386	4	2	2	2342	2343	
0	2389	4	2	2	2344	2345	
0	2392	4	2	2	2346	2347	
0	2395	4	2	2	2348	2349	
0	2398	4	3	2	7897	7191	
0	2402	4	1	2	7893	7899	
0	2403	4	1	2	7900	7224	
0	2404	4	2	2	7826	7901	
0	2407	4	2	2	2357	2358	
0	2410	4	3	2	7287	7902	
0	2414	4	3	2	7904	6807	
0	2418	4	3	2	7906	6839	
0	2422	4	3	2	7908	6871	
0	2426	4	3	2	7910	6903	
0	2430	4	3	2	7912	6935	
0	2434	4	3	2	7914	6967	
0	2438	4	3	2	7916	6999	
0	2442	4	3	2	7918	7031	
0	2446	4	3	2	7920	7063	
0	2450	4	3	2	7922	7095	
0	2454	4	3	2	7924	7127	
0	2458	4	3	2	7926	7159	
0	2462	4	1	2	7898	7928	
0	2463	4	1	2	7929	7192	
0	2464	4	2	2	7853	7930	
0	2467	4	2	2	2402	2403	
0	2470	4	3	2	7933	7931	
0	2474	4	1	2	7288	7935	
0	2475	4	1	2	7936	7903	
0	2476	4	1	2	7905	7938	
0	2477	4	1	2	7939	6808	
0	2478	4	2	2	7858	7940	
0	2481	4	1	2	7907	7941	
0	2482	4	1	2	7942	6840	
0	2483	4	2	2	7861	7943	
0	2486	4	1	2	7909	7944	
0	2487	4	1	2	7945	6872	
0	2488	4	2	2	7864	7946	
0	2491	4	1	2	7911	7947	
0	2492	4	1	2	7948	6904	
0	2493	4	2	2	7867	7949	
0	2496	4	1	2	7913	7950	
0	2497	4	1	2	7951	6936	
0	2498	4	2	2	7870	7952	
0	2501	4	1	2	7915	7953	
0	2502	4	1	2	7954	6968	
0	2503	4	2	2	7873	7955	
0	2506	4	1	2	7917	7956	
0	2507	4	1	2	7957	7000	
0	2508	4	2	2	7876	7958	
0	2511	4	1	2	7919	7959	
0	2512	4	1	2	7960	7032	
0	2513	4	2	2	7879	7961	
0	2516	4	1	2	7921	7962	
0	2517	4	1	2	7963	7064	
0	2518	4	2	2	7882	7964	
0	2521	4	1	2	7923	7965	
0	2522	4	1	2	7966	7096	
0	2523	4	2	2	7885	7967	
0	2526	4	1	2	7925	7968	
0	2527	4	1	2	7969	7128	
0	2528	4	2	2	7888	7970	
0	2531	4	1	2	7927	7971	
0	2532	4	1	2	7972	7160	
0	2533	4	2	2	7891	7973	
0	2536	4	2	2	2462	2463	
0	2539	4	3	2	7976	7974	
0	2543	4	1	2	7934	7978	
0	2544	4	1	2	7979	7932	
0	2545	4	2	2	2474	2475	
3	2548	4	0	2	2476	2477	
0	2549	4	2	2	2481	2482	
0	2552	4	2	2	2486	2487	
0	2555	4	2	2	2491	2492	
0	2558	4	2	2	2496	2497	
0	2561	4	2	2	2501	2502	
0	2564	4	2	2	2506	2507	
0	2567	4	2	2	2511	2512	
0	2570	4	2	2	2516	2517	
0	2573	4	2	2	2521	2522	
0	2576	4	2	2	2526	2527	
0	2579	4	2	2	2531	2532	
0	2582	4	3	2	8005	8003	
0	2586	4	1	2	7977	8007	
0	2587	4	1	2	8008	7975	
0	2588	4	2	2	2543	2544	
0	2591	4	3	2	8010	7257	
0	2595	4	3	2	8012	7981	
0	2599	4	3	2	8014	7983	
0	2603	4	3	2	8016	7985	
0	2607	4	3	2	8018	7987	
0	2611	4	3	2	8020	7989	
0	2615	4	3	2	8022	7991	
0	2619	4	3	2	8024	7993	
0	2623	4	3	2	8026	7995	
0	2627	4	3	2	8028	7997	
0	2631	4	3	2	8030	7999	
0	2635	4	3	2	8032	8001	
0	2639	4	1	2	8006	8034	
0	2640	4	1	2	8035	8004	
0	2641	4	2	2	2586	2587	
0	2644	4	3	2	8037	7225	
0	2648	4	1	2	8011	8039	
0	2649	4	1	2	8040	7258	
0	2650	4	2	2	7937	8041	
0	2653	4	1	2	8013	8042	
0	2654	4	1	2	8043	7982	
0	2655	4	1	2	8015	8045	
0	2656	4	1	2	8046	7984	
0	2657	4	1	2	8017	8048	
0	2658	4	1	2	8049	7986	
0	2659	4	1	2	8019	8051	
0	2660	4	1	2	8052	7988	
0	2661	4	1	2	8021	8054	
0	2662	4	1	2	8055	7990	
0	2663	4	1	2	8023	8057	
0	2664	4	1	2	8058	7992	
0	2665	4	1	2	8025	8060	
0	2666	4	1	2	8061	7994	
0	2667	4	1	2	8027	8063	
0	2668	4	1	2	8064	7996	
0	2669	4	1	2	8029	8066	
0	2670	4	1	2	8067	7998	
0	2671	4	1	2	8031	8069	
0	2672	4	1	2	8070	8000	
0	2673	4	1	2	8033	8072	
0	2674	4	1	2	8073	8002	
0	2675	4	2	2	2639	2640	
0	2678	4	3	2	8075	7193	
0	2682	4	1	2	8038	8077	
0	2683	4	1	2	8078	7226	
0	2684	4	2	2	7980	8079	
0	2687	4	2	2	2648	2649	
0	2690	4	3	2	7289	8080	
0	2694	4	2	2	2653	2654	
0	2697	4	2	2	2655	2656	
0	2700	4	2	2	2657	2658	
0	2703	4	2	2	2659	2660	
0	2706	4	2	2	2661	2662	
0	2709	4	2	2	2663	2664	
0	2712	4	2	2	2665	2666	
0	2715	4	2	2	2667	2668	
0	2718	4	2	2	2669	2670	
0	2721	4	2	2	2671	2672	
0	2724	4	2	2	2673	2674	
0	2727	4	3	2	8082	7161	
0	2731	4	1	2	8076	8084	
0	2732	4	1	2	8085	7194	
0	2733	4	2	2	8009	8086	
0	2736	4	2	2	2682	2683	
0	2739	4	3	2	8089	8087	
0	2743	4	1	2	7290	8091	
0	2744	4	1	2	8092	8081	
0	2745	4	3	2	8094	6809	
0	2749	4	3	2	8096	6841	
0	2753	4	3	2	8098	6873	
0	2757	4	3	2	8100	6905	
0	2761	4	3	2	8102	6937	
0	2765	4	3	2	8104	6969	
0	2769	4	3	2	8106	7001	
0	2773	4	3	2	8108	7033	
0	2777	4	3	2	8110	7065	
0	2781	4	3	2	8112	7097	
0	2785	4	3	2	8114	7129	
0	2789	4	1	2	8083	8116	
0	2790	4	1	2	8117	7162	
0	2791	4	2	2	8036	8118	
0	2794	4	2	2	2731	2732	
0	2797	4	3	2	8121	8119	
0	2801	4	1	2	8090	8123	
0	2802	4	1	2	8124	8088	
0	2803	4	2	2	2743	2744	
0	2806	4	1	2	8095	8126	
0	2807	4	1	2	8127	6810	
0	2808	4	2	2	8044	8128	
0	2811	4	1	2	8097	8129	
0	2812	4	1	2	8130	6842	
0	2813	4	2	2	8047	8131	
0	2816	4	1	2	8099	8132	
0	2817	4	1	2	8133	6874	
0	2818	4	2	2	8050	8134	
0	2821	4	1	2	8101	8135	
0	2822	4	1	2	8136	6906	
0	2823	4	2	2	8053	8137	
0	2826	4	1	2	8103	8138	
0	2827	4	1	2	8139	6938	
0	2828	4	2	2	8056	8140	
0	2831	4	1	2	8105	8141	
0	2832	4	1	2	8142	6970	
0	2833	4	2	2	8059	8143	
0	2836	4	1	2	8107	8144	
0	2837	4	1	2	8145	7002	
0	2838	4	2	2	8062	8146	
0	2841	4	1	2	8109	8147	
0	2842	4	1	2	8148	7034	
0	2843	4	2	2	8065	8149	
0	2846	4	1	2	8111	8150	
0	2847	4	1	2	8151	7066	
0	2848	4	2	2	8068	8152	
0	2851	4	1	2	8113	8153	
0	2852	4	1	2	8154	7098	
0	2853	4	2	2	8071	8155	
0	2856	4	1	2	8115	8156	
0	2857	4	1	2	8157	7130	
0	2858	4	2	2	8074	8158	
0	2861	4	2	2	2789	2790	
0	2864	4	3	2	8161	8159	
0	2868	4	1	2	8122	8163	
0	2869	4	1	2	8164	8120	
0	2870	4	2	2	2801	2802	
0	2873	4	3	2	8166	7259	
3	2877	4	0	2	2806	2807	
0	2878	4	2	2	2811	2812	
0	2881	4	2	2	2816	2817	
0	2884	4	2	2	2821	2822	
0	2887	4	2	2	2826	2827	
0	2890	4	2	2	2831	2832	
0	2893	4	2	2	2836	2837	
0	2896	4	2	2	2841	2842	
0	2899	4	2	2	2846	2847	
0	2902	4	2	2	2851	2852	
0	2905	4	2	2	2856	2857	
0	2908	4	3	2	8190	8188	
0	2912	4	1	2	8162	8192	
0	2913	4	1	2	8193	8160	
0	2914	4	2	2	2868	2869	
0	2917	4	3	2	8195	7227	
0	2921	4	1	2	8167	8197	
0	2922	4	1	2	8198	7260	
0	2923	4	2	2	8093	8199	
0	2926	4	3	2	8200	8168	
0	2930	4	3	2	8202	8170	
0	2934	4	3	2	8204	8172	
0	2938	4	3	2	8206	8174	
0	2942	4	3	2	8208	8176	
0	2946	4	3	2	8210	8178	
0	2950	4	3	2	8212	8180	
0	2954	4	3	2	8214	8182	
0	2958	4	3	2	8216	8184	
0	2962	4	3	2	8218	8186	
0	2966	4	1	2	8191	8220	
0	2967	4	1	2	8221	8189	
0	2968	4	2	2	2912	2913	
0	2971	4	3	2	8223	7195	
0	2975	4	1	2	8196	8225	
0	2976	4	1	2	8226	7228	
0	2977	4	2	2	8125	8227	
0	2980	4	2	2	2921	2922	
0	2983	4	3	2	7291	8228	
0	2987	4	1	2	8201	8230	
0	2988	4	1	2	8231	8169	
0	2989	4	1	2	8203	8233	
0	2990	4	1	2	8234	8171	
0	2991	4	1	2	8205	8236	
0	2992	4	1	2	8237	8173	
0	2993	4	1	2	8207	8239	
0	2994	4	1	2	8240	8175	
0	2995	4	1	2	8209	8242	
0	2996	4	1	2	8243	8177	
0	2997	4	1	2	8211	8245	
0	2998	4	1	2	8246	8179	
0	2999	4	1	2	8213	8248	
0	3000	4	1	2	8249	8181	
0	3001	4	1	2	8215	8251	
0	3002	4	1	2	8252	8183	
0	3003	4	1	2	8217	8254	
0	3004	4	1	2	8255	8185	
0	3005	4	1	2	8219	8257	
0	3006	4	1	2	8258	8187	
0	3007	4	2	2	2966	2967	
0	3010	4	3	2	8260	7163	
0	3014	4	1	2	8224	8262	
0	3015	4	1	2	8263	7196	
0	3016	4	2	2	8165	8264	
0	3019	4	2	2	2975	2976	
0	3022	4	3	2	8267	8265	
0	3026	4	1	2	7292	8269	
0	3027	4	1	2	8270	8229	
0	3028	4	2	2	2987	2988	
0	3031	4	2	2	2989	2990	
0	3034	4	2	2	2991	2992	
0	3037	4	2	2	2993	2994	
0	3040	4	2	2	2995	2996	
0	3043	4	2	2	2997	2998	
0	3046	4	2	2	2999	3000	
0	3049	4	2	2	3001	3002	
0	3052	4	2	2	3003	3004	
0	3055	4	2	2	3005	3006	
0	3058	4	3	2	8272	7131	
0	3062	4	1	2	8261	8274	
0	3063	4	1	2	8275	7164	
0	3064	4	2	2	8194	8276	
0	3067	4	2	2	3014	3015	
0	3070	4	3	2	8279	8277	
0	3074	4	1	2	8268	8281	
0	3075	4	1	2	8282	8266	
0	3076	4	2	2	3026	3027	
0	3079	4	3	2	8284	6811	
0	3083	4	3	2	8286	6843	
0	3087	4	3	2	8288	6875	
0	3091	4	3	2	8290	6907	
0	3095	4	3	2	8292	6939	
0	3099	4	3	2	8294	6971	
0	3103	4	3	2	8296	7003	
0	3107	4	3	2	8298	7035	
0	3111	4	3	2	8300	7067	
0	3115	4	3	2	8302	7099	
0	3119	4	1	2	8273	8304	
0	3120	4	1	2	8305	7132	
0	3121	4	2	2	8222	8306	
0	3124	4	2	2	3062	3063	
0	3127	4	3	2	8309	8307	
0	3131	4	1	2	8280	8311	
0	3132	4	1	2	8312	8278	
0	3133	4	2	2	3074	3075	
0	3136	4	3	2	8314	7261	
0	3140	4	1	2	8285	8316	
0	3141	4	1	2	8317	6812	
0	3142	4	2	2	8232	8318	
0	3145	4	1	2	8287	8319	
0	3146	4	1	2	8320	6844	
0	3147	4	2	2	8235	8321	
0	3150	4	1	2	8289	8322	
0	3151	4	1	2	8323	6876	
0	3152	4	2	2	8238	8324	
0	3155	4	1	2	8291	8325	
0	3156	4	1	2	8326	6908	
0	3157	4	2	2	8241	8327	
0	3160	4	1	2	8293	8328	
0	3161	4	1	2	8329	6940	
0	3162	4	2	2	8244	8330	
0	3165	4	1	2	8295	8331	
0	3166	4	1	2	8332	6972	
0	3167	4	2	2	8247	8333	
0	3170	4	1	2	8297	8334	
0	3171	4	1	2	8335	7004	
0	3172	4	2	2	8250	8336	
0	3175	4	1	2	8299	8337	
0	3176	4	1	2	8338	7036	
0	3177	4	2	2	8253	8339	
0	3180	4	1	2	8301	8340	
0	3181	4	1	2	8341	7068	
0	3182	4	2	2	8256	8342	
0	3185	4	1	2	8303	8343	
0	3186	4	1	2	8344	7100	
0	3187	4	2	2	8259	8345	
0	3190	4	2	2	3119	3120	
0	3193	4	3	2	8348	8346	
0	3197	4	1	2	8310	8350	
0	3198	4	1	2	8351	8308	
0	3199	4	2	2	3131	3132	
0	3202	4	3	2	8353	7229	
0	3206	4	1	2	8315	8355	
0	3207	4	1	2	8356	7262	
0	3208	4	2	2	8271	8357	
3	3211	4	0	2	3140	3141	
0	3212	4	2	2	3145	3146	
0	3215	4	2	2	3150	3151	
0	3218	4	2	2	3155	3156	
0	3221	4	2	2	3160	3161	
0	3224	4	2	2	3165	3166	
0	3227	4	2	2	3170	3171	
0	3230	4	2	2	3175	3176	
0	3233	4	2	2	3180	3181	
0	3236	4	2	2	3185	3186	
0	3239	4	3	2	8378	8376	
0	3243	4	1	2	8349	8380	
0	3244	4	1	2	8381	8347	
0	3245	4	2	2	3197	3198	
0	3248	4	3	2	8383	7197	
0	3252	4	1	2	8354	8385	
0	3253	4	1	2	8386	7230	
0	3254	4	2	2	8283	8387	
0	3257	4	2	2	3206	3207	
0	3260	4	3	2	7293	8388	
0	3264	4	3	2	8390	8358	
0	3268	4	3	2	8392	8360	
0	3272	4	3	2	8394	8362	
0	3276	4	3	2	8396	8364	
0	3280	4	3	2	8398	8366	
0	3284	4	3	2	8400	8368	
0	3288	4	3	2	8402	8370	
0	3292	4	3	2	8404	8372	
0	3296	4	3	2	8406	8374	
0	3300	4	1	2	8379	8408	
0	3301	4	1	2	8409	8377	
0	3302	4	2	2	3243	3244	
0	3305	4	3	2	8411	7165	
0	3309	4	1	2	8384	8413	
0	3310	4	1	2	8414	7198	
0	3311	4	2	2	8313	8415	
0	3314	4	2	2	3252	3253	
0	3317	4	3	2	8418	8416	
0	3321	4	1	2	7294	8420	
0	3322	4	1	2	8421	8389	
0	3323	4	1	2	8391	8423	
0	3324	4	1	2	8424	8359	
0	3325	4	1	2	8393	8426	
0	3326	4	1	2	8427	8361	
0	3327	4	1	2	8395	8429	
0	3328	4	1	2	8430	8363	
0	3329	4	1	2	8397	8432	
0	3330	4	1	2	8433	8365	
0	3331	4	1	2	8399	8435	
0	3332	4	1	2	8436	8367	
0	3333	4	1	2	8401	8438	
0	3334	4	1	2	8439	8369	
0	3335	4	1	2	8403	8441	
0	3336	4	1	2	8442	8371	
0	3337	4	1	2	8405	8444	
0	3338	4	1	2	8445	8373	
0	3339	4	1	2	8407	8447	
0	3340	4	1	2	8448	8375	
0	3341	4	2	2	3300	3301	
0	3344	4	3	2	8450	7133	
0	3348	4	1	2	8412	8452	
0	3349	4	1	2	8453	7166	
0	3350	4	2	2	8352	8454	
0	3353	4	2	2	3309	3310	
0	3356	4	3	2	8457	8455	
0	3360	4	1	2	8419	8459	
0	3361	4	1	2	8460	8417	
0	3362	4	2	2	3321	3322	
0	3365	4	2	2	3323	3324	
0	3368	4	2	2	3325	3326	
0	3371	4	2	2	3327	3328	
0	3374	4	2	2	3329	3330	
0	3377	4	2	2	3331	3332	
0	3380	4	2	2	3333	3334	
0	3383	4	2	2	3335	3336	
0	3386	4	2	2	3337	3338	
0	3389	4	2	2	3339	3340	
0	3392	4	3	2	8462	7101	
0	3396	4	1	2	8451	8464	
0	3397	4	1	2	8465	7134	
0	3398	4	2	2	8382	8466	
0	3401	4	2	2	3348	3349	
0	3404	4	3	2	8469	8467	
0	3408	4	1	2	8458	8471	
0	3409	4	1	2	8472	8456	
0	3410	4	2	2	3360	3361	
0	3413	4	3	2	8474	7263	
0	3417	4	3	2	8476	6813	
0	3421	4	3	2	8478	6845	
0	3425	4	3	2	8480	6877	
0	3429	4	3	2	8482	6909	
0	3433	4	3	2	8484	6941	
0	3437	4	3	2	8486	6973	
0	3441	4	3	2	8488	7005	
0	3445	4	3	2	8490	7037	
0	3449	4	3	2	8492	7069	
0	3453	4	1	2	8463	8494	
0	3454	4	1	2	8495	7102	
0	3455	4	2	2	8410	8496	
0	3458	4	2	2	3396	3397	
0	3461	4	3	2	8499	8497	
0	3465	4	1	2	8470	8501	
0	3466	4	1	2	8502	8468	
0	3467	4	2	2	3408	3409	
0	3470	4	3	2	8504	7231	
0	3474	4	1	2	8475	8506	
0	3475	4	1	2	8507	7264	
0	3476	4	2	2	8422	8508	
0	3479	4	1	2	8477	8509	
0	3480	4	1	2	8510	6814	
0	3481	4	2	2	8425	8511	
0	3484	4	1	2	8479	8512	
0	3485	4	1	2	8513	6846	
0	3486	4	2	2	8428	8514	
0	3489	4	1	2	8481	8515	
0	3490	4	1	2	8516	6878	
0	3491	4	2	2	8431	8517	
0	3494	4	1	2	8483	8518	
0	3495	4	1	2	8519	6910	
0	3496	4	2	2	8434	8520	
0	3499	4	1	2	8485	8521	
0	3500	4	1	2	8522	6942	
0	3501	4	2	2	8437	8523	
0	3504	4	1	2	8487	8524	
0	3505	4	1	2	8525	6974	
0	3506	4	2	2	8440	8526	
0	3509	4	1	2	8489	8527	
0	3510	4	1	2	8528	7006	
0	3511	4	2	2	8443	8529	
0	3514	4	1	2	8491	8530	
0	3515	4	1	2	8531	7038	
0	3516	4	2	2	8446	8532	
0	3519	4	1	2	8493	8533	
0	3520	4	1	2	8534	7070	
0	3521	4	2	2	8449	8535	
0	3524	4	2	2	3453	3454	
0	3527	4	3	2	8538	8536	
0	3531	4	1	2	8500	8540	
0	3532	4	1	2	8541	8498	
0	3533	4	2	2	3465	3466	
0	3536	4	3	2	8543	7199	
0	3540	4	1	2	8505	8545	
0	3541	4	1	2	8546	7232	
0	3542	4	2	2	8461	8547	
0	3545	4	2	2	3474	3475	
0	3548	4	3	2	7295	8548	
3	3552	4	0	2	3479	3480	
0	3553	4	2	2	3484	3485	
0	3556	4	2	2	3489	3490	
0	3559	4	2	2	3494	3495	
0	3562	4	2	2	3499	3500	
0	3565	4	2	2	3504	3505	
0	3568	4	2	2	3509	3510	
0	3571	4	2	2	3514	3515	
0	3574	4	2	2	3519	3520	
0	3577	4	3	2	8568	8566	
0	3581	4	1	2	8539	8570	
0	3582	4	1	2	8571	8537	
0	3583	4	2	2	3531	3532	
0	3586	4	3	2	8573	7167	
0	3590	4	1	2	8544	8575	
0	3591	4	1	2	8576	7200	
0	3592	4	2	2	8473	8577	
0	3595	4	2	2	3540	3541	
0	3598	4	3	2	8580	8578	
0	3602	4	1	2	7296	8582	
0	3603	4	1	2	8583	8549	
0	3604	4	3	2	8585	8550	
0	3608	4	3	2	8587	8552	
0	3612	4	3	2	8589	8554	
0	3616	4	3	2	8591	8556	
0	3620	4	3	2	8593	8558	
0	3624	4	3	2	8595	8560	
0	3628	4	3	2	8597	8562	
0	3632	4	3	2	8599	8564	
0	3636	4	1	2	8569	8601	
0	3637	4	1	2	8602	8567	
0	3638	4	2	2	3581	3582	
0	3641	4	3	2	8604	7135	
0	3645	4	1	2	8574	8606	
0	3646	4	1	2	8607	7168	
0	3647	4	2	2	8503	8608	
0	3650	4	2	2	3590	3591	
0	3653	4	3	2	8611	8609	
0	3657	4	1	2	8581	8613	
0	3658	4	1	2	8614	8579	
0	3659	4	2	2	3602	3603	
0	3662	4	1	2	8586	8616	
0	3663	4	1	2	8617	8551	
0	3664	4	1	2	8588	8619	
0	3665	4	1	2	8620	8553	
0	3666	4	1	2	8590	8622	
0	3667	4	1	2	8623	8555	
0	3668	4	1	2	8592	8625	
0	3669	4	1	2	8626	8557	
0	3670	4	1	2	8594	8628	
0	3671	4	1	2	8629	8559	
0	3672	4	1	2	8596	8631	
0	3673	4	1	2	8632	8561	
0	3674	4	1	2	8598	8634	
0	3675	4	1	2	8635	8563	
0	3676	4	1	2	8600	8637	
0	3677	4	1	2	8638	8565	
0	3678	4	2	2	3636	3637	
0	3681	4	3	2	8640	7103	
0	3685	4	1	2	8605	8642	
0	3686	4	1	2	8643	7136	
0	3687	4	2	2	8542	8644	
0	3690	4	2	2	3645	3646	
0	3693	4	3	2	8647	8645	
0	3697	4	1	2	8612	8649	
0	3698	4	1	2	8650	8610	
0	3699	4	2	2	3657	3658	
0	3702	4	3	2	8652	7265	
0	3706	4	2	2	3662	3663	
0	3709	4	2	2	3664	3665	
0	3712	4	2	2	3666	3667	
0	3715	4	2	2	3668	3669	
0	3718	4	2	2	3670	3671	
0	3721	4	2	2	3672	3673	
0	3724	4	2	2	3674	3675	
0	3727	4	2	2	3676	3677	
0	3730	4	3	2	8654	7071	
0	3734	4	1	2	8641	8656	
0	3735	4	1	2	8657	7104	
0	3736	4	2	2	8572	8658	
0	3739	4	2	2	3685	3686	
0	3742	4	3	2	8661	8659	
0	3746	4	1	2	8648	8663	
0	3747	4	1	2	8664	8646	
0	3748	4	2	2	3697	3698	
0	3751	4	3	2	8666	7233	
0	3755	4	1	2	8653	8668	
0	3756	4	1	2	8669	7266	
0	3757	4	2	2	8584	8670	
0	3760	4	3	2	8671	6815	
0	3764	4	3	2	8673	6847	
0	3768	4	3	2	8675	6879	
0	3772	4	3	2	8677	6911	
0	3776	4	3	2	8679	6943	
0	3780	4	3	2	8681	6975	
0	3784	4	3	2	8683	7007	
0	3788	4	3	2	8685	7039	
0	3792	4	1	2	8655	8687	
0	3793	4	1	2	8688	7072	
0	3794	4	2	2	8603	8689	
0	3797	4	2	2	3734	3735	
0	3800	4	3	2	8692	8690	
0	3804	4	1	2	8662	8694	
0	3805	4	1	2	8695	8660	
0	3806	4	2	2	3746	3747	
0	3809	4	3	2	8697	7201	
0	3813	4	1	2	8667	8699	
0	3814	4	1	2	8700	7234	
0	3815	4	2	2	8615	8701	
0	3818	4	2	2	3755	3756	
0	3821	4	3	2	7297	8702	
0	3825	4	1	2	8672	8704	
0	3826	4	1	2	8705	6816	
0	3827	4	2	2	8618	8706	
0	3830	4	1	2	8674	8707	
0	3831	4	1	2	8708	6848	
0	3832	4	2	2	8621	8709	
0	3835	4	1	2	8676	8710	
0	3836	4	1	2	8711	6880	
0	3837	4	2	2	8624	8712	
0	3840	4	1	2	8678	8713	
0	3841	4	1	2	8714	6912	
0	3842	4	2	2	8627	8715	
0	3845	4	1	2	8680	8716	
0	3846	4	1	2	8717	6944	
0	3847	4	2	2	8630	8718	
0	3850	4	1	2	8682	8719	
0	3851	4	1	2	8720	6976	
0	3852	4	2	2	8633	8721	
0	3855	4	1	2	8684	8722	
0	3856	4	1	2	8723	7008	
0	3857	4	2	2	8636	8724	
0	3860	4	1	2	8686	8725	
0	3861	4	1	2	8726	7040	
0	3862	4	2	2	8639	8727	
0	3865	4	2	2	3792	3793	
0	3868	4	3	2	8730	8728	
0	3872	4	1	2	8693	8732	
0	3873	4	1	2	8733	8691	
0	3874	4	2	2	3804	3805	
0	3877	4	3	2	8735	7169	
0	3881	4	1	2	8698	8737	
0	3882	4	1	2	8738	7202	
0	3883	4	2	2	8651	8739	
0	3886	4	2	2	3813	3814	
0	3889	4	3	2	8742	8740	
0	3893	4	1	2	7298	8744	
0	3894	4	1	2	8745	8703	
3	3895	4	0	2	3825	3826	
0	3896	4	2	2	3830	3831	
0	3899	4	2	2	3835	3836	
0	3902	4	2	2	3840	3841	
0	3905	4	2	2	3845	3846	
0	3908	4	2	2	3850	3851	
0	3911	4	2	2	3855	3856	
0	3914	4	2	2	3860	3861	
0	3917	4	3	2	8763	8761	
0	3921	4	1	2	8731	8765	
0	3922	4	1	2	8766	8729	
0	3923	4	2	2	3872	3873	
0	3926	4	3	2	8768	7137	
0	3930	4	1	2	8736	8770	
0	3931	4	1	2	8771	7170	
0	3932	4	2	2	8665	8772	
0	3935	4	2	2	3881	3882	
0	3938	4	3	2	8775	8773	
0	3942	4	1	2	8743	8777	
0	3943	4	1	2	8778	8741	
0	3944	4	2	2	3893	3894	
0	3947	4	3	2	8780	8747	
0	3951	4	3	2	8782	8749	
0	3955	4	3	2	8784	8751	
0	3959	4	3	2	8786	8753	
0	3963	4	3	2	8788	8755	
0	3967	4	3	2	8790	8757	
0	3971	4	3	2	8792	8759	
0	3975	4	1	2	8764	8794	
0	3976	4	1	2	8795	8762	
0	3977	4	2	2	3921	3922	
0	3980	4	3	2	8797	7105	
0	3984	4	1	2	8769	8799	
0	3985	4	1	2	8800	7138	
0	3986	4	2	2	8696	8801	
0	3989	4	2	2	3930	3931	
0	3992	4	3	2	8804	8802	
0	3996	4	1	2	8776	8806	
0	3997	4	1	2	8807	8774	
0	3998	4	2	2	3942	3943	
0	4001	4	3	2	8809	7267	
0	4005	4	1	2	8781	8811	
0	4006	4	1	2	8812	8748	
0	4007	4	1	2	8783	8814	
0	4008	4	1	2	8815	8750	
0	4009	4	1	2	8785	8817	
0	4010	4	1	2	8818	8752	
0	4011	4	1	2	8787	8820	
0	4012	4	1	2	8821	8754	
0	4013	4	1	2	8789	8823	
0	4014	4	1	2	8824	8756	
0	4015	4	1	2	8791	8826	
0	4016	4	1	2	8827	8758	
0	4017	4	1	2	8793	8829	
0	4018	4	1	2	8830	8760	
0	4019	4	2	2	3975	3976	
0	4022	4	3	2	8832	7073	
0	4026	4	1	2	8798	8834	
0	4027	4	1	2	8835	7106	
0	4028	4	2	2	8734	8836	
0	4031	4	2	2	3984	3985	
0	4034	4	3	2	8839	8837	
0	4038	4	1	2	8805	8841	
0	4039	4	1	2	8842	8803	
0	4040	4	2	2	3996	3997	
0	4043	4	3	2	8844	7235	
0	4047	4	1	2	8810	8846	
0	4048	4	1	2	8847	7268	
0	4049	4	2	2	8746	8848	
0	4052	4	2	2	4005	4006	
0	4055	4	2	2	4007	4008	
0	4058	4	2	2	4009	4010	
0	4061	4	2	2	4011	4012	
0	4064	4	2	2	4013	4014	
0	4067	4	2	2	4015	4016	
0	4070	4	2	2	4017	4018	
0	4073	4	3	2	8849	7041	
0	4077	4	1	2	8833	8851	
0	4078	4	1	2	8852	7074	
0	4079	4	2	2	8767	8853	
0	4082	4	2	2	4026	4027	
0	4085	4	3	2	8856	8854	
0	4089	4	1	2	8840	8858	
0	4090	4	1	2	8859	8838	
0	4091	4	2	2	4038	4039	
0	4094	4	3	2	8861	7203	
0	4098	4	1	2	8845	8863	
0	4099	4	1	2	8864	7236	
0	4100	4	2	2	8779	8865	
0	4103	4	2	2	4047	4048	
0	4106	4	3	2	7299	8866	
0	4110	4	3	2	8868	6817	
0	4114	4	3	2	8870	6849	
0	4118	4	3	2	8872	6881	
0	4122	4	3	2	8874	6913	
0	4126	4	3	2	8876	6945	
0	4130	4	3	2	8878	6977	
0	4134	4	3	2	8880	7009	
0	4138	4	1	2	8850	8882	
0	4139	4	1	2	8883	7042	
0	4140	4	2	2	8796	8884	
0	4143	4	2	2	4077	4078	
0	4146	4	3	2	8887	8885	
0	4150	4	1	2	8857	8889	
0	4151	4	1	2	8890	8855	
0	4152	4	2	2	4089	4090	
0	4155	4	3	2	8892	7171	
0	4159	4	1	2	8862	8894	
0	4160	4	1	2	8895	7204	
0	4161	4	2	2	8808	8896	
0	4164	4	2	2	4098	4099	
0	4167	4	3	2	8899	8897	
0	4171	4	1	2	7300	8901	
0	4172	4	1	2	8902	8867	
0	4173	4	1	2	8869	8904	
0	4174	4	1	2	8905	6818	
0	4175	4	2	2	8813	8906	
0	4178	4	1	2	8871	8907	
0	4179	4	1	2	8908	6850	
0	4180	4	2	2	8816	8909	
0	4183	4	1	2	8873	8910	
0	4184	4	1	2	8911	6882	
0	4185	4	2	2	8819	8912	
0	4188	4	1	2	8875	8913	
0	4189	4	1	2	8914	6914	
0	4190	4	2	2	8822	8915	
0	4193	4	1	2	8877	8916	
0	4194	4	1	2	8917	6946	
0	4195	4	2	2	8825	8918	
0	4198	4	1	2	8879	8919	
0	4199	4	1	2	8920	6978	
0	4200	4	2	2	8828	8921	
0	4203	4	1	2	8881	8922	
0	4204	4	1	2	8923	7010	
0	4205	4	2	2	8831	8924	
0	4208	4	2	2	4138	4139	
0	4211	4	3	2	8927	8925	
0	4215	4	1	2	8888	8929	
0	4216	4	1	2	8930	8886	
0	4217	4	2	2	4150	4151	
0	4220	4	3	2	8932	7139	
0	4224	4	1	2	8893	8934	
0	4225	4	1	2	8935	7172	
0	4226	4	2	2	8843	8936	
0	4229	4	2	2	4159	4160	
0	4232	4	3	2	8939	8937	
0	4236	4	1	2	8900	8941	
0	4237	4	1	2	8942	8898	
0	4238	4	2	2	4171	4172	
3	4241	4	0	2	4173	4174	
0	4242	4	2	2	4178	4179	
0	4245	4	2	2	4183	4184	
0	4248	4	2	2	4188	4189	
0	4251	4	2	2	4193	4194	
0	4254	4	2	2	4198	4199	
0	4257	4	2	2	4203	4204	
0	4260	4	3	2	8958	8956	
0	4264	4	1	2	8928	8960	
0	4265	4	1	2	8961	8926	
0	4266	4	2	2	4215	4216	
0	4269	4	3	2	8963	7107	
0	4273	4	1	2	8933	8965	
0	4274	4	1	2	8966	7140	
0	4275	4	2	2	8860	8967	
0	4278	4	2	2	4224	4225	
0	4281	4	3	2	8970	8968	
0	4285	4	1	2	8940	8972	
0	4286	4	1	2	8973	8938	
0	4287	4	2	2	4236	4237	
0	4290	4	3	2	8975	7269	
0	4294	4	3	2	8977	8944	
0	4298	4	3	2	8979	8946	
0	4302	4	3	2	8981	8948	
0	4306	4	3	2	8983	8950	
0	4310	4	3	2	8985	8952	
0	4314	4	3	2	8987	8954	
0	4318	4	1	2	8959	8989	
0	4319	4	1	2	8990	8957	
0	4320	4	2	2	4264	4265	
0	4323	4	3	2	8992	7075	
0	4327	4	1	2	8964	8994	
0	4328	4	1	2	8995	7108	
0	4329	4	2	2	8891	8996	
0	4332	4	2	2	4273	4274	
0	4335	4	3	2	8999	8997	
0	4339	4	1	2	8971	9001	
0	4340	4	1	2	9002	8969	
0	4341	4	2	2	4285	4286	
0	4344	4	3	2	9004	7237	
0	4348	4	1	2	8976	9006	
0	4349	4	1	2	9007	7270	
0	4350	4	2	2	8903	9008	
0	4353	4	1	2	8978	9009	
0	4354	4	1	2	9010	8945	
0	4355	4	1	2	8980	9012	
0	4356	4	1	2	9013	8947	
0	4357	4	1	2	8982	9015	
0	4358	4	1	2	9016	8949	
0	4359	4	1	2	8984	9018	
0	4360	4	1	2	9019	8951	
0	4361	4	1	2	8986	9021	
0	4362	4	1	2	9022	8953	
0	4363	4	1	2	8988	9024	
0	4364	4	1	2	9025	8955	
0	4365	4	2	2	4318	4319	
0	4368	4	3	2	9027	7043	
0	4372	4	1	2	8993	9029	
0	4373	4	1	2	9030	7076	
0	4374	4	2	2	8931	9031	
0	4377	4	2	2	4327	4328	
0	4380	4	3	2	9034	9032	
0	4384	4	1	2	9000	9036	
0	4385	4	1	2	9037	8998	
0	4386	4	2	2	4339	4340	
0	4389	4	3	2	9039	7205	
0	4393	4	1	2	9005	9041	
0	4394	4	1	2	9042	7238	
0	4395	4	2	2	8943	9043	
0	4398	4	2	2	4348	4349	
0	4401	4	3	2	7301	9044	
0	4405	4	2	2	4353	4354	
0	4408	4	2	2	4355	4356	
0	4411	4	2	2	4357	4358	
0	4414	4	2	2	4359	4360	
0	4417	4	2	2	4361	4362	
0	4420	4	2	2	4363	4364	
0	4423	4	3	2	9046	7011	
0	4427	4	1	2	9028	9048	
0	4428	4	1	2	9049	7044	
0	4429	4	2	2	8962	9050	
0	4432	4	2	2	4372	4373	
0	4435	4	3	2	9053	9051	
0	4439	4	1	2	9035	9055	
0	4440	4	1	2	9056	9033	
0	4441	4	2	2	4384	4385	
0	4444	4	3	2	9058	7173	
0	4448	4	1	2	9040	9060	
0	4449	4	1	2	9061	7206	
0	4450	4	2	2	8974	9062	
0	4453	4	2	2	4393	4394	
0	4456	4	3	2	9065	9063	
0	4460	4	1	2	7302	9067	
0	4461	4	1	2	9068	9045	
0	4462	4	3	2	9070	6819	
0	4466	4	3	2	9072	6851	
0	4470	4	3	2	9074	6883	
0	4474	4	3	2	9076	6915	
0	4478	4	3	2	9078	6947	
0	4482	4	3	2	9080	6979	
0	4486	4	1	2	9047	9082	
0	4487	4	1	2	9083	7012	
0	4488	4	2	2	8991	9084	
0	4491	4	2	2	4427	4428	
0	4494	4	3	2	9087	9085	
0	4498	4	1	2	9054	9089	
0	4499	4	1	2	9090	9052	
0	4500	4	2	2	4439	4440	
0	4503	4	3	2	9092	7141	
0	4507	4	1	2	9059	9094	
0	4508	4	1	2	9095	7174	
0	4509	4	2	2	9003	9096	
0	4512	4	2	2	4448	4449	
0	4515	4	3	2	9099	9097	
0	4519	4	1	2	9066	9101	
0	4520	4	1	2	9102	9064	
0	4521	4	2	2	4460	4461	
0	4524	4	1	2	9071	9104	
0	4525	4	1	2	9105	6820	
0	4526	4	2	2	9011	9106	
0	4529	4	1	2	9073	9107	
0	4530	4	1	2	9108	6852	
0	4531	4	2	2	9014	9109	
0	4534	4	1	2	9075	9110	
0	4535	4	1	2	9111	6884	
0	4536	4	2	2	9017	9112	
0	4539	4	1	2	9077	9113	
0	4540	4	1	2	9114	6916	
0	4541	4	2	2	9020	9115	
0	4544	4	1	2	9079	9116	
0	4545	4	1	2	9117	6948	
0	4546	4	2	2	9023	9118	
0	4549	4	1	2	9081	9119	
0	4550	4	1	2	9120	6980	
0	4551	4	2	2	9026	9121	
0	4554	4	2	2	4486	4487	
0	4557	4	3	2	9124	9122	
0	4561	4	1	2	9088	9126	
0	4562	4	1	2	9127	9086	
0	4563	4	2	2	4498	4499	
0	4566	4	3	2	9129	7109	
0	4570	4	1	2	9093	9131	
0	4571	4	1	2	9132	7142	
0	4572	4	2	2	9038	9133	
0	4575	4	2	2	4507	4508	
0	4578	4	3	2	9136	9134	
0	4582	4	1	2	9100	9138	
0	4583	4	1	2	9139	9098	
0	4584	4	2	2	4519	4520	
0	4587	4	3	2	9141	7271	
3	4591	4	0	2	4524	4525	
0	4592	4	2	2	4529	4530	
0	4595	4	2	2	4534	4535	
0	4598	4	2	2	4539	4540	
0	4601	4	2	2	4544	4545	
0	4604	4	2	2	4549	4550	
0	4607	4	3	2	9155	9153	
0	4611	4	1	2	9125	9157	
0	4612	4	1	2	9158	9123	
0	4613	4	2	2	4561	4562	
0	4616	4	3	2	9160	7077	
0	4620	4	1	2	9130	9162	
0	4621	4	1	2	9163	7110	
0	4622	4	2	2	9057	9164	
0	4625	4	2	2	4570	4571	
0	4628	4	3	2	9167	9165	
0	4632	4	1	2	9137	9169	
0	4633	4	1	2	9170	9135	
0	4634	4	2	2	4582	4583	
0	4637	4	3	2	9172	7239	
0	4641	4	1	2	9142	9174	
0	4642	4	1	2	9175	7272	
0	4643	4	2	2	9069	9176	
0	4646	4	3	2	9177	9143	
0	4650	4	3	2	9179	9145	
0	4654	4	3	2	9181	9147	
0	4658	4	3	2	9183	9149	
0	4662	4	3	2	9185	9151	
0	4666	4	1	2	9156	9187	
0	4667	4	1	2	9188	9154	
0	4668	4	2	2	4611	4612	
0	4671	4	3	2	9190	7045	
0	4675	4	1	2	9161	9192	
0	4676	4	1	2	9193	7078	
0	4677	4	2	2	9091	9194	
0	4680	4	2	2	4620	4621	
0	4683	4	3	2	9197	9195	
0	4687	4	1	2	9168	9199	
0	4688	4	1	2	9200	9166	
0	4689	4	2	2	4632	4633	
0	4692	4	3	2	9202	7207	
0	4696	4	1	2	9173	9204	
0	4697	4	1	2	9205	7240	
0	4698	4	2	2	9103	9206	
0	4701	4	2	2	4641	4642	
0	4704	4	3	2	7303	9207	
0	4708	4	1	2	9178	9209	
0	4709	4	1	2	9210	9144	
0	4710	4	1	2	9180	9212	
0	4711	4	1	2	9213	9146	
0	4712	4	1	2	9182	9215	
0	4713	4	1	2	9216	9148	
0	4714	4	1	2	9184	9218	
0	4715	4	1	2	9219	9150	
0	4716	4	1	2	9186	9221	
0	4717	4	1	2	9222	9152	
0	4718	4	2	2	4666	4667	
0	4721	4	3	2	9224	7013	
0	4725	4	1	2	9191	9226	
0	4726	4	1	2	9227	7046	
0	4727	4	2	2	9128	9228	
0	4730	4	2	2	4675	4676	
0	4733	4	3	2	9231	9229	
0	4737	4	1	2	9198	9233	
0	4738	4	1	2	9234	9196	
0	4739	4	2	2	4687	4688	
0	4742	4	3	2	9236	7175	
0	4746	4	1	2	9203	9238	
0	4747	4	1	2	9239	7208	
0	4748	4	2	2	9140	9240	
0	4751	4	2	2	4696	4697	
0	4754	4	3	2	9243	9241	
0	4758	4	1	2	7304	9245	
0	4759	4	1	2	9246	9208	
0	4760	4	2	2	4708	4709	
0	4763	4	2	2	4710	4711	
0	4766	4	2	2	4712	4713	
0	4769	4	2	2	4714	4715	
0	4772	4	2	2	4716	4717	
0	4775	4	3	2	9248	6981	
0	4779	4	1	2	9225	9250	
0	4780	4	1	2	9251	7014	
0	4781	4	2	2	9159	9252	
0	4784	4	2	2	4725	4726	
0	4787	4	3	2	9255	9253	
0	4791	4	1	2	9232	9257	
0	4792	4	1	2	9258	9230	
0	4793	4	2	2	4737	4738	
0	4796	4	3	2	9260	7143	
0	4800	4	1	2	9237	9262	
0	4801	4	1	2	9263	7176	
0	4802	4	2	2	9171	9264	
0	4805	4	2	2	4746	4747	
0	4808	4	3	2	9267	9265	
0	4812	4	1	2	9244	9269	
0	4813	4	1	2	9270	9242	
0	4814	4	2	2	4758	4759	
0	4817	4	3	2	9272	6821	
0	4821	4	3	2	9274	6853	
0	4825	4	3	2	9276	6885	
0	4829	4	3	2	9278	6917	
0	4833	4	3	2	9280	6949	
0	4837	4	1	2	9249	9282	
0	4838	4	1	2	9283	6982	
0	4839	4	2	2	9189	9284	
0	4842	4	2	2	4779	4780	
0	4845	4	3	2	9287	9285	
0	4849	4	1	2	9256	9289	
0	4850	4	1	2	9290	9254	
0	4851	4	2	2	4791	4792	
0	4854	4	3	2	9292	7111	
0	4858	4	1	2	9261	9294	
0	4859	4	1	2	9295	7144	
0	4860	4	2	2	9201	9296	
0	4863	4	2	2	4800	4801	
0	4866	4	3	2	9299	9297	
0	4870	4	1	2	9268	9301	
0	4871	4	1	2	9302	9266	
0	4872	4	2	2	4812	4813	
0	4875	4	3	2	9304	7273	
0	4879	4	1	2	9273	9306	
0	4880	4	1	2	9307	6822	
0	4881	4	2	2	9211	9308	
0	4884	4	1	2	9275	9309	
0	4885	4	1	2	9310	6854	
0	4886	4	2	2	9214	9311	
0	4889	4	1	2	9277	9312	
0	4890	4	1	2	9313	6886	
0	4891	4	2	2	9217	9314	
0	4894	4	1	2	9279	9315	
0	4895	4	1	2	9316	6918	
0	4896	4	2	2	9220	9317	
0	4899	4	1	2	9281	9318	
0	4900	4	1	2	9319	6950	
0	4901	4	2	2	9223	9320	
0	4904	4	2	2	4837	4838	
0	4907	4	3	2	9323	9321	
0	4911	4	1	2	9288	9325	
0	4912	4	1	2	9326	9286	
0	4913	4	2	2	4849	4850	
0	4916	4	3	2	9328	7079	
0	4920	4	1	2	9293	9330	
0	4921	4	1	2	9331	7112	
0	4922	4	2	2	9235	9332	
0	4925	4	2	2	4858	4859	
0	4928	4	3	2	9335	9333	
0	4932	4	1	2	9300	9337	
0	4933	4	1	2	9338	9298	
0	4934	4	2	2	4870	4871	
0	4937	4	3	2	9340	7241	
0	4941	4	1	2	9305	9342	
0	4942	4	1	2	9343	7274	
0	4943	4	2	2	9247	9344	
3	4946	4	0	2	4879	4880	
0	4947	4	2	2	4884	4885	
0	4950	4	2	2	4889	4890	
0	4953	4	2	2	4894	4895	
0	4956	4	2	2	4899	4900	
0	4959	4	3	2	9355	9353	
0	4963	4	1	2	9324	9357	
0	4964	4	1	2	9358	9322	
0	4965	4	2	2	4911	4912	
0	4968	4	3	2	9360	7047	
0	4972	4	1	2	9329	9362	
0	4973	4	1	2	9363	7080	
0	4974	4	2	2	9259	9364	
0	4977	4	2	2	4920	4921	
0	4980	4	3	2	9367	9365	
0	4984	4	1	2	9336	9369	
0	4985	4	1	2	9370	9334	
0	4986	4	2	2	4932	4933	
0	4989	4	3	2	9372	7209	
0	4993	4	1	2	9341	9374	
0	4994	4	1	2	9375	7242	
0	4995	4	2	2	9271	9376	
0	4998	4	2	2	4941	4942	
0	5001	4	3	2	7305	9377	
0	5005	4	3	2	9379	9345	
0	5009	4	3	2	9381	9347	
0	5013	4	3	2	9383	9349	
0	5017	4	3	2	9385	9351	
0	5021	4	1	2	9356	9387	
0	5022	4	1	2	9388	9354	
0	5023	4	2	2	4963	4964	
0	5026	4	3	2	9390	7015	
0	5030	4	1	2	9361	9392	
0	5031	4	1	2	9393	7048	
0	5032	4	2	2	9291	9394	
0	5035	4	2	2	4972	4973	
0	5038	4	3	2	9397	9395	
0	5042	4	1	2	9368	9399	
0	5043	4	1	2	9400	9366	
0	5044	4	2	2	4984	4985	
0	5047	4	3	2	9402	7177	
0	5051	4	1	2	9373	9404	
0	5052	4	1	2	9405	7210	
0	5053	4	2	2	9303	9406	
0	5056	4	2	2	4993	4994	
0	5059	4	3	2	9409	9407	
0	5063	4	1	2	7306	9411	
0	5064	4	1	2	9412	9378	
0	5065	4	1	2	9380	9414	
0	5066	4	1	2	9415	9346	
0	5067	4	1	2	9382	9417	
0	5068	4	1	2	9418	9348	
0	5069	4	1	2	9384	9420	
0	5070	4	1	2	9421	9350	
0	5071	4	1	2	9386	9423	
0	5072	4	1	2	9424	9352	
0	5073	4	2	2	5021	5022	
0	5076	4	3	2	9426	6983	
0	5080	4	1	2	9391	9428	
0	5081	4	1	2	9429	7016	
0	5082	4	2	2	9327	9430	
0	5085	4	2	2	5030	5031	
0	5088	4	3	2	9433	9431	
0	5092	4	1	2	9398	9435	
0	5093	4	1	2	9436	9396	
0	5094	4	2	2	5042	5043	
0	5097	4	3	2	9438	7145	
0	5101	4	1	2	9403	9440	
0	5102	4	1	2	9441	7178	
0	5103	4	2	2	9339	9442	
0	5106	4	2	2	5051	5052	
0	5109	4	3	2	9445	9443	
0	5113	4	1	2	9410	9447	
0	5114	4	1	2	9448	9408	
0	5115	4	2	2	5063	5064	
0	5118	4	2	2	5065	5066	
0	5121	4	2	2	5067	5068	
0	5124	4	2	2	5069	5070	
0	5127	4	2	2	5071	5072	
0	5130	4	3	2	9450	6951	
0	5134	4	1	2	9427	9452	
0	5135	4	1	2	9453	6984	
0	5136	4	2	2	9359	9454	
0	5139	4	2	2	5080	5081	
0	5142	4	3	2	9457	9455	
0	5146	4	1	2	9434	9459	
0	5147	4	1	2	9460	9432	
0	5148	4	2	2	5092	5093	
0	5151	4	3	2	9462	7113	
0	5155	4	1	2	9439	9464	
0	5156	4	1	2	9465	7146	
0	5157	4	2	2	9371	9466	
0	5160	4	2	2	5101	5102	
0	5163	4	3	2	9469	9467	
0	5167	4	1	2	9446	9471	
0	5168	4	1	2	9472	9444	
0	5169	4	2	2	5113	5114	
0	5172	4	3	2	9474	7275	
0	5176	4	3	2	9476	6823	
0	5180	4	3	2	9478	6855	
0	5184	4	3	2	9480	6887	
0	5188	4	3	2	9482	6919	
0	5192	4	1	2	9451	9484	
0	5193	4	1	2	9485	6952	
0	5194	4	2	2	9389	9486	
0	5197	4	2	2	5134	5135	
0	5200	4	3	2	9489	9487	
0	5204	4	1	2	9458	9491	
0	5205	4	1	2	9492	9456	
0	5206	4	2	2	5146	5147	
0	5209	4	3	2	9494	7081	
0	5213	4	1	2	9463	9496	
0	5214	4	1	2	9497	7114	
0	5215	4	2	2	9401	9498	
0	5218	4	2	2	5155	5156	
0	5221	4	3	2	9501	9499	
0	5225	4	1	2	9470	9503	
0	5226	4	1	2	9504	9468	
0	5227	4	2	2	5167	5168	
0	5230	4	3	2	9506	7243	
0	5234	4	1	2	9475	9508	
0	5235	4	1	2	9509	7276	
0	5236	4	2	2	9413	9510	
0	5239	4	1	2	9477	9511	
0	5240	4	1	2	9512	6824	
0	5241	4	2	2	9416	9513	
0	5244	4	1	2	9479	9514	
0	5245	4	1	2	9515	6856	
0	5246	4	2	2	9419	9516	
0	5249	4	1	2	9481	9517	
0	5250	4	1	2	9518	6888	
0	5251	4	2	2	9422	9519	
0	5254	4	1	2	9483	9520	
0	5255	4	1	2	9521	6920	
0	5256	4	2	2	9425	9522	
0	5259	4	2	2	5192	5193	
0	5262	4	3	2	9525	9523	
0	5266	4	1	2	9490	9527	
0	5267	4	1	2	9528	9488	
0	5268	4	2	2	5204	5205	
0	5271	4	3	2	9530	7049	
0	5275	4	1	2	9495	9532	
0	5276	4	1	2	9533	7082	
0	5277	4	2	2	9437	9534	
0	5280	4	2	2	5213	5214	
0	5283	4	3	2	9537	9535	
0	5287	4	1	2	9502	9539	
0	5288	4	1	2	9540	9500	
0	5289	4	2	2	5225	5226	
0	5292	4	3	2	9542	7211	
0	5296	4	1	2	9507	9544	
0	5297	4	1	2	9545	7244	
0	5298	4	2	2	9449	9546	
0	5301	4	2	2	5234	5235	
0	5304	4	3	2	7307	9547	
3	5308	4	0	2	5239	5240	
0	5309	4	2	2	5244	5245	
0	5312	4	2	2	5249	5250	
0	5315	4	2	2	5254	5255	
0	5318	4	3	2	9557	9555	
0	5322	4	1	2	9526	9559	
0	5323	4	1	2	9560	9524	
0	5324	4	2	2	5266	5267	
0	5327	4	3	2	9562	7017	
0	5331	4	1	2	9531	9564	
0	5332	4	1	2	9565	7050	
0	5333	4	2	2	9461	9566	
0	5336	4	2	2	5275	5276	
0	5339	4	3	2	9569	9567	
0	5343	4	1	2	9538	9571	
0	5344	4	1	2	9572	9536	
0	5345	4	2	2	5287	5288	
0	5348	4	3	2	9574	7179	
0	5352	4	1	2	9543	9576	
0	5353	4	1	2	9577	7212	
0	5354	4	2	2	9473	9578	
0	5357	4	2	2	5296	5297	
0	5360	4	3	2	9581	9579	
0	5364	4	1	2	7308	9583	
0	5365	4	1	2	9584	9548	
0	5366	4	3	2	9586	9549	
0	5370	4	3	2	9588	9551	
0	5374	4	3	2	9590	9553	
0	5378	4	1	2	9558	9592	
0	5379	4	1	2	9593	9556	
0	5380	4	2	2	5322	5323	
0	5383	4	3	2	9595	6985	
0	5387	4	1	2	9563	9597	
0	5388	4	1	2	9598	7018	
0	5389	4	2	2	9493	9599	
0	5392	4	2	2	5331	5332	
0	5395	4	3	2	9602	9600	
0	5399	4	1	2	9570	9604	
0	5400	4	1	2	9605	9568	
0	5401	4	2	2	5343	5344	
0	5404	4	3	2	9607	7147	
0	5408	4	1	2	9575	9609	
0	5409	4	1	2	9610	7180	
0	5410	4	2	2	9505	9611	
0	5413	4	2	2	5352	5353	
0	5416	4	3	2	9614	9612	
0	5420	4	1	2	9582	9616	
0	5421	4	1	2	9617	9580	
0	5422	4	2	2	5364	5365	
0	5425	4	1	2	9587	9619	
0	5426	4	1	2	9620	9550	
0	5427	4	1	2	9589	9622	
0	5428	4	1	2	9623	9552	
0	5429	4	1	2	9591	9625	
0	5430	4	1	2	9626	9554	
0	5431	4	2	2	5378	5379	
0	5434	4	3	2	9628	6953	
0	5438	4	1	2	9596	9630	
0	5439	4	1	2	9631	6986	
0	5440	4	2	2	9529	9632	
0	5443	4	2	2	5387	5388	
0	5446	4	3	2	9635	9633	
0	5450	4	1	2	9603	9637	
0	5451	4	1	2	9638	9601	
0	5452	4	2	2	5399	5400	
0	5455	4	3	2	9640	7115	
0	5459	4	1	2	9608	9642	
0	5460	4	1	2	9643	7148	
0	5461	4	2	2	9541	9644	
0	5464	4	2	2	5408	5409	
0	5467	4	3	2	9647	9645	
0	5471	4	1	2	9615	9649	
0	5472	4	1	2	9650	9613	
0	5473	4	2	2	5420	5421	
0	5476	4	3	2	9652	7277	
0	5480	4	2	2	5425	5426	
0	5483	4	2	2	5427	5428	
0	5486	4	2	2	5429	5430	
0	5489	4	3	2	9654	6921	
0	5493	4	1	2	9629	9656	
0	5494	4	1	2	9657	6954	
0	5495	4	2	2	9561	9658	
0	5498	4	2	2	5438	5439	
0	5501	4	3	2	9661	9659	
0	5505	4	1	2	9636	9663	
0	5506	4	1	2	9664	9634	
0	5507	4	2	2	5450	5451	
0	5510	4	3	2	9666	7083	
0	5514	4	1	2	9641	9668	
0	5515	4	1	2	9669	7116	
0	5516	4	2	2	9573	9670	
0	5519	4	2	2	5459	5460	
0	5522	4	3	2	9673	9671	
0	5526	4	1	2	9648	9675	
0	5527	4	1	2	9676	9646	
0	5528	4	2	2	5471	5472	
0	5531	4	3	2	9678	7245	
0	5535	4	1	2	9653	9680	
0	5536	4	1	2	9681	7278	
0	5537	4	2	2	9585	9682	
0	5540	4	3	2	9683	6825	
0	5544	4	3	2	9685	6857	
0	5548	4	3	2	9687	6889	
0	5552	4	1	2	9655	9689	
0	5553	4	1	2	9690	6922	
0	5554	4	2	2	9594	9691	
0	5557	4	2	2	5493	5494	
0	5560	4	3	2	9694	9692	
0	5564	4	1	2	9662	9696	
0	5565	4	1	2	9697	9660	
0	5566	4	2	2	5505	5506	
0	5569	4	3	2	9699	7051	
0	5573	4	1	2	9667	9701	
0	5574	4	1	2	9702	7084	
0	5575	4	2	2	9606	9703	
0	5578	4	2	2	5514	5515	
0	5581	4	3	2	9706	9704	
0	5585	4	1	2	9674	9708	
0	5586	4	1	2	9709	9672	
0	5587	4	2	2	5526	5527	
0	5590	4	3	2	9711	7213	
0	5594	4	1	2	9679	9713	
0	5595	4	1	2	9714	7246	
0	5596	4	2	2	9618	9715	
0	5599	4	2	2	5535	5536	
0	5602	4	3	2	7309	9716	
0	5606	4	1	2	9684	9718	
0	5607	4	1	2	9719	6826	
0	5608	4	2	2	9621	9720	
0	5611	4	1	2	9686	9721	
0	5612	4	1	2	9722	6858	
0	5613	4	2	2	9624	9723	
0	5616	4	1	2	9688	9724	
0	5617	4	1	2	9725	6890	
0	5618	4	2	2	9627	9726	
0	5621	4	2	2	5552	5553	
0	5624	4	3	2	9729	9727	
0	5628	4	1	2	9695	9731	
0	5629	4	1	2	9732	9693	
0	5630	4	2	2	5564	5565	
0	5633	4	3	2	9734	7019	
0	5637	4	1	2	9700	9736	
0	5638	4	1	2	9737	7052	
0	5639	4	2	2	9639	9738	
0	5642	4	2	2	5573	5574	
0	5645	4	3	2	9741	9739	
0	5649	4	1	2	9707	9743	
0	5650	4	1	2	9744	9705	
0	5651	4	2	2	5585	5586	
0	5654	4	3	2	9746	7181	
0	5658	4	1	2	9712	9748	
0	5659	4	1	2	9749	7214	
0	5660	4	2	2	9651	9750	
0	5663	4	2	2	5594	5595	
0	5666	4	3	2	9753	9751	
0	5670	4	1	2	7310	9755	
0	5671	4	1	2	9756	9717	
3	5672	4	0	2	5606	5607	
0	5673	4	2	2	5611	5612	
0	5676	4	2	2	5616	5617	
0	5679	4	3	2	9764	9762	
0	5683	4	1	2	9730	9766	
0	5684	4	1	2	9767	9728	
0	5685	4	2	2	5628	5629	
0	5688	4	3	2	9769	6987	
0	5692	4	1	2	9735	9771	
0	5693	4	1	2	9772	7020	
0	5694	4	2	2	9665	9773	
0	5697	4	2	2	5637	5638	
0	5700	4	3	2	9776	9774	
0	5704	4	1	2	9742	9778	
0	5705	4	1	2	9779	9740	
0	5706	4	2	2	5649	5650	
0	5709	4	3	2	9781	7149	
0	5713	4	1	2	9747	9783	
0	5714	4	1	2	9784	7182	
0	5715	4	2	2	9677	9785	
0	5718	4	2	2	5658	5659	
0	5721	4	3	2	9788	9786	
0	5725	4	1	2	9754	9790	
0	5726	4	1	2	9791	9752	
0	5727	4	2	2	5670	5671	
0	5730	4	3	2	9793	9758	
0	5734	4	3	2	9795	9760	
0	5738	4	1	2	9765	9797	
0	5739	4	1	2	9798	9763	
0	5740	4	2	2	5683	5684	
0	5743	4	3	2	9800	6955	
0	5747	4	1	2	9770	9802	
0	5748	4	1	2	9803	6988	
0	5749	4	2	2	9698	9804	
0	5752	4	2	2	5692	5693	
0	5755	4	3	2	9807	9805	
0	5759	4	1	2	9777	9809	
0	5760	4	1	2	9810	9775	
0	5761	4	2	2	5704	5705	
0	5764	4	3	2	9812	7117	
0	5768	4	1	2	9782	9814	
0	5769	4	1	2	9815	7150	
0	5770	4	2	2	9710	9816	
0	5773	4	2	2	5713	5714	
0	5776	4	3	2	9819	9817	
0	5780	4	1	2	9789	9821	
0	5781	4	1	2	9822	9787	
0	5782	4	2	2	5725	5726	
0	5785	4	1	2	9794	9826	
0	5786	4	1	2	9827	9759	
0	5787	4	1	2	9796	9829	
0	5788	4	1	2	9830	9761	
0	5789	4	2	2	5738	5739	
0	5792	4	3	2	9832	6923	
0	5796	4	1	2	9801	9834	
0	5797	4	1	2	9835	6956	
0	5798	4	2	2	9733	9836	
0	5801	4	2	2	5747	5748	
0	5804	4	3	2	9839	9837	
0	5808	4	1	2	9808	9841	
0	5809	4	1	2	9842	9806	
0	5810	4	2	2	5759	5760	
0	5813	4	3	2	9844	7085	
0	5817	4	1	2	9813	9846	
0	5818	4	1	2	9847	7118	
0	5819	4	2	2	9745	9848	
0	5822	4	2	2	5768	5769	
0	5825	4	3	2	9851	9849	
0	5829	4	1	2	9820	9853	
0	5830	4	1	2	9854	9818	
0	5831	4	2	2	5780	5781	
0	5834	4	2	2	5785	5786	
0	5837	4	2	2	5787	5788	
0	5840	4	3	2	9858	6891	
0	5844	4	1	2	9833	9860	
0	5845	4	1	2	9861	6924	
0	5846	4	2	2	9768	9862	
0	5849	4	2	2	5796	5797	
0	5852	4	3	2	9865	9863	
0	5856	4	1	2	9840	9867	
0	5857	4	1	2	9868	9838	
0	5858	4	2	2	5808	5809	
0	5861	4	3	2	9870	7053	
0	5865	4	1	2	9845	9872	
0	5866	4	1	2	9873	7086	
0	5867	4	2	2	9780	9874	
0	5870	4	2	2	5817	5818	
0	5873	4	3	2	9877	9875	
0	5877	4	1	2	9852	9879	
0	5878	4	1	2	9880	9850	
0	5879	4	2	2	5829	5830	
0	5882	4	3	2	9884	6827	
0	5886	4	3	2	9886	6859	
0	5890	4	1	2	9859	9888	
0	5891	4	1	2	9889	6892	
0	5892	4	2	2	9799	9890	
0	5895	4	2	2	5844	5845	
0	5898	4	3	2	9893	9891	
0	5902	4	1	2	9866	9895	
0	5903	4	1	2	9896	9864	
0	5904	4	2	2	5856	5857	
0	5907	4	3	2	9898	7021	
0	5911	4	1	2	9871	9900	
0	5912	4	1	2	9901	7054	
0	5913	4	2	2	9811	9902	
0	5916	4	2	2	5865	5866	
0	5919	4	3	2	9905	9903	
0	5923	4	1	2	9878	9907	
0	5924	4	1	2	9908	9876	
0	5925	4	2	2	5877	5878	
0	5928	4	1	2	9885	9912	
0	5929	4	1	2	9913	6828	
0	5930	4	2	2	9828	9914	
0	5933	4	1	2	9887	9915	
0	5934	4	1	2	9916	6860	
0	5935	4	2	2	9831	9917	
0	5938	4	2	2	5890	5891	
0	5941	4	3	2	9920	9918	
0	5945	4	1	2	9894	9922	
0	5946	4	1	2	9923	9892	
0	5947	4	2	2	5902	5903	
0	5950	4	3	2	9925	6989	
0	5954	4	1	2	9899	9927	
0	5955	4	1	2	9928	7022	
0	5956	4	2	2	9843	9929	
0	5959	4	2	2	5911	5912	
0	5962	4	3	2	9932	9930	
0	5966	4	1	2	9906	9934	
0	5967	4	1	2	9935	9904	
0	5968	4	2	2	5923	5924	
3	5971	4	0	2	5928	5929	
0	5972	4	2	2	5933	5934	
0	5975	4	3	2	9943	9941	
0	5979	4	1	2	9921	9945	
0	5980	4	1	2	9946	9919	
0	5981	4	2	2	5945	5946	
0	5984	4	3	2	9948	6957	
0	5988	4	1	2	9926	9950	
0	5989	4	1	2	9951	6990	
0	5990	4	2	2	9869	9952	
0	5993	4	2	2	5954	5955	
0	5996	4	3	2	9955	9953	
0	6000	4	1	2	9933	9957	
0	6001	4	1	2	9958	9931	
0	6002	4	2	2	5966	5967	
0	6005	4	3	2	9962	9939	
0	6009	4	1	2	9944	9964	
0	6010	4	1	2	9965	9942	
0	6011	4	2	2	5979	5980	
0	6014	4	3	2	9967	6925	
0	6018	4	1	2	9949	9969	
0	6019	4	1	2	9970	6958	
0	6020	4	2	2	9897	9971	
0	6023	4	2	2	5988	5989	
0	6026	4	3	2	9974	9972	
0	6030	4	1	2	9956	9976	
0	6031	4	1	2	9977	9954	
0	6032	4	2	2	6000	6001	
0	6035	4	1	2	9963	9981	
0	6036	4	1	2	9982	9940	
0	6037	4	2	2	6009	6010	
0	6040	4	3	2	9984	6893	
0	6044	4	1	2	9968	9986	
0	6045	4	1	2	9987	6926	
0	6046	4	2	2	9924	9988	
0	6049	4	2	2	6018	6019	
0	6052	4	3	2	9991	9989	
0	6056	4	1	2	9975	9993	
0	6057	4	1	2	9994	9973	
0	6058	4	2	2	6030	6031	
0	6061	4	2	2	6035	6036	
0	6064	4	3	2	9998	6861	
0	6068	4	1	2	9985	10000	
0	6069	4	1	2	10001	6894	
0	6070	4	2	2	9947	10002	
0	6073	4	2	2	6044	6045	
0	6076	4	3	2	10005	10003	
0	6080	4	1	2	9992	10007	
0	6081	4	1	2	10008	9990	
0	6082	4	2	2	6056	6057	
0	6085	4	3	2	10012	6829	
0	6089	4	1	2	9999	10014	
0	6090	4	1	2	10015	6862	
0	6091	4	2	2	9966	10016	
0	6094	4	2	2	6068	6069	
0	6097	4	3	2	10019	10017	
0	6101	4	1	2	10006	10021	
0	6102	4	1	2	10022	10004	
0	6103	4	2	2	6080	6081	
0	6106	4	1	2	10013	10026	
0	6107	4	1	2	10027	6830	
0	6108	4	2	2	9983	10028	
0	6111	4	2	2	6089	6090	
0	6114	4	3	2	10031	10029	
0	6118	4	1	2	10020	10033	
0	6119	4	1	2	10034	10018	
0	6120	4	2	2	6101	6102	
3	6123	4	0	2	6106	6107	
0	6124	4	3	2	10040	10038	
0	6128	4	1	2	10032	10042	
0	6129	4	1	2	10043	10030	
0	6130	4	2	2	6118	6119	
0	6133	4	1	2	10041	10047	
0	6134	4	1	2	10048	10039	
0	6135	4	2	2	6128	6129	
0	6138	4	2	2	6133	6134	
0	6141	5	3	1	10054	
0	6145	4	1	2	10055	10056	
0	6146	5	1	1	10057	
0	6147	4	2	2	10049	10058	
3	6150	4	0	2	6145	6146	
0	6151	4	3	2	10052	10059	
0	6155	4	1	2	10053	10061	
0	6156	4	1	2	10062	10060	
0	6157	4	2	2	10044	10063	
3	6160	4	0	2	6155	6156	
0	6161	4	3	2	10050	10064	
0	6165	4	1	2	10051	10066	
0	6166	4	1	2	10067	10065	
0	6167	4	2	2	10035	10068	
3	6170	4	0	2	6165	6166	
0	6171	4	3	2	10045	10069	
0	6175	4	1	2	10046	10071	
0	6176	4	1	2	10072	10070	
0	6177	4	2	2	10023	10073	
3	6180	4	0	2	6175	6176	
0	6181	4	3	2	10036	10074	
0	6185	4	1	2	10037	10076	
0	6186	4	1	2	10077	10075	
0	6187	4	2	2	10009	10078	
3	6190	4	0	2	6185	6186	
0	6191	4	3	2	10024	10079	
0	6195	4	1	2	10025	10081	
0	6196	4	1	2	10082	10080	
0	6197	4	2	2	9995	10083	
3	6200	4	0	2	6195	6196	
0	6201	4	3	2	10010	10084	
0	6205	4	1	2	10011	10086	
0	6206	4	1	2	10087	10085	
0	6207	4	2	2	9978	10088	
3	6210	4	0	2	6205	6206	
0	6211	4	3	2	9996	10089	
0	6215	4	1	2	9997	10091	
0	6216	4	1	2	10092	10090	
0	6217	4	2	2	9959	10093	
3	6220	4	0	2	6215	6216	
0	6221	4	3	2	9979	10094	
0	6225	4	1	2	9980	10096	
0	6226	4	1	2	10097	10095	
0	6227	4	2	2	9936	10098	
3	6230	4	0	2	6225	6226	
0	6231	4	3	2	9960	10099	
0	6235	4	1	2	9961	10101	
0	6236	4	1	2	10102	10100	
0	6237	4	2	2	9909	10103	
3	6240	4	0	2	6235	6236	
0	6241	4	3	2	9937	10104	
0	6245	4	1	2	9938	10106	
0	6246	4	1	2	10107	10105	
0	6247	4	2	2	9881	10108	
3	6250	4	0	2	6245	6246	
0	6251	4	3	2	9910	10109	
0	6255	4	1	2	9911	10111	
0	6256	4	1	2	10112	10110	
0	6257	4	2	2	9855	10113	
3	6260	4	0	2	6255	6256	
0	6261	4	3	2	9882	10114	
0	6265	4	1	2	9883	10116	
0	6266	4	1	2	10117	10115	
0	6267	4	2	2	9823	10118	
3	6270	4	0	2	6265	6266	
0	6271	4	3	2	9856	10119	
0	6275	4	1	2	9857	10121	
0	6276	4	1	2	10122	10120	
0	6277	4	2	2	9792	10123	
3	6280	4	0	2	6275	6276	
0	6281	4	3	2	9824	10124	
0	6285	4	1	2	9825	10126	
0	6286	4	1	2	10127	10125	
3	6287	4	0	2	9757	10128	
3	6288	4	0	2	6285	6286	
2	6289	1	1			
2	6290	1	1			
2	6291	1	1			
2	6292	1	1			
2	6293	1	1			
2	6294	1	1			
2	6295	1	1			
2	6296	1	1			
2	6297	1	1			
2	6298	1	1			
2	6299	1	1			
2	6300	1	1			
2	6301	1	1			
2	6302	1	1			
2	6303	1	1			
2	6304	1	1			
2	6305	1	18			
2	6306	1	18			
2	6307	1	18			
2	6308	1	18			
2	6309	1	18			
2	6310	1	18			
2	6311	1	18			
2	6312	1	18			
2	6313	1	18			
2	6314	1	18			
2	6315	1	18			
2	6316	1	18			
2	6317	1	18			
2	6318	1	18			
2	6319	1	18			
2	6320	1	18			
2	6321	1	35			
2	6322	1	35			
2	6323	1	35			
2	6324	1	35			
2	6325	1	35			
2	6326	1	35			
2	6327	1	35			
2	6328	1	35			
2	6329	1	35			
2	6330	1	35			
2	6331	1	35			
2	6332	1	35			
2	6333	1	35			
2	6334	1	35			
2	6335	1	35			
2	6336	1	35			
2	6337	1	52			
2	6338	1	52			
2	6339	1	52			
2	6340	1	52			
2	6341	1	52			
2	6342	1	52			
2	6343	1	52			
2	6344	1	52			
2	6345	1	52			
2	6346	1	52			
2	6347	1	52			
2	6348	1	52			
2	6349	1	52			
2	6350	1	52			
2	6351	1	52			
2	6352	1	52			
2	6353	1	69			
2	6354	1	69			
2	6355	1	69			
2	6356	1	69			
2	6357	1	69			
2	6358	1	69			
2	6359	1	69			
2	6360	1	69			
2	6361	1	69			
2	6362	1	69			
2	6363	1	69			
2	6364	1	69			
2	6365	1	69			
2	6366	1	69			
2	6367	1	69			
2	6368	1	69			
2	6369	1	86			
2	6370	1	86			
2	6371	1	86			
2	6372	1	86			
2	6373	1	86			
2	6374	1	86			
2	6375	1	86			
2	6376	1	86			
2	6377	1	86			
2	6378	1	86			
2	6379	1	86			
2	6380	1	86			
2	6381	1	86			
2	6382	1	86			
2	6383	1	86			
2	6384	1	86			
2	6385	1	103			
2	6386	1	103			
2	6387	1	103			
2	6388	1	103			
2	6389	1	103			
2	6390	1	103			
2	6391	1	103			
2	6392	1	103			
2	6393	1	103			
2	6394	1	103			
2	6395	1	103			
2	6396	1	103			
2	6397	1	103			
2	6398	1	103			
2	6399	1	103			
2	6400	1	103			
2	6401	1	120			
2	6402	1	120			
2	6403	1	120			
2	6404	1	120			
2	6405	1	120			
2	6406	1	120			
2	6407	1	120			
2	6408	1	120			
2	6409	1	120			
2	6410	1	120			
2	6411	1	120			
2	6412	1	120			
2	6413	1	120			
2	6414	1	120			
2	6415	1	120			
2	6416	1	120			
2	6417	1	137			
2	6418	1	137			
2	6419	1	137			
2	6420	1	137			
2	6421	1	137			
2	6422	1	137			
2	6423	1	137			
2	6424	1	137			
2	6425	1	137			
2	6426	1	137			
2	6427	1	137			
2	6428	1	137			
2	6429	1	137			
2	6430	1	137			
2	6431	1	137			
2	6432	1	137			
2	6433	1	154			
2	6434	1	154			
2	6435	1	154			
2	6436	1	154			
2	6437	1	154			
2	6438	1	154			
2	6439	1	154			
2	6440	1	154			
2	6441	1	154			
2	6442	1	154			
2	6443	1	154			
2	6444	1	154			
2	6445	1	154			
2	6446	1	154			
2	6447	1	154			
2	6448	1	154			
2	6449	1	171			
2	6450	1	171			
2	6451	1	171			
2	6452	1	171			
2	6453	1	171			
2	6454	1	171			
2	6455	1	171			
2	6456	1	171			
2	6457	1	171			
2	6458	1	171			
2	6459	1	171			
2	6460	1	171			
2	6461	1	171			
2	6462	1	171			
2	6463	1	171			
2	6464	1	171			
2	6465	1	188			
2	6466	1	188			
2	6467	1	188			
2	6468	1	188			
2	6469	1	188			
2	6470	1	188			
2	6471	1	188			
2	6472	1	188			
2	6473	1	188			
2	6474	1	188			
2	6475	1	188			
2	6476	1	188			
2	6477	1	188			
2	6478	1	188			
2	6479	1	188			
2	6480	1	188			
2	6481	1	205			
2	6482	1	205			
2	6483	1	205			
2	6484	1	205			
2	6485	1	205			
2	6486	1	205			
2	6487	1	205			
2	6488	1	205			
2	6489	1	205			
2	6490	1	205			
2	6491	1	205			
2	6492	1	205			
2	6493	1	205			
2	6494	1	205			
2	6495	1	205			
2	6496	1	205			
2	6497	1	222			
2	6498	1	222			
2	6499	1	222			
2	6500	1	222			
2	6501	1	222			
2	6502	1	222			
2	6503	1	222			
2	6504	1	222			
2	6505	1	222			
2	6506	1	222			
2	6507	1	222			
2	6508	1	222			
2	6509	1	222			
2	6510	1	222			
2	6511	1	222			
2	6512	1	222			
2	6513	1	239			
2	6514	1	239			
2	6515	1	239			
2	6516	1	239			
2	6517	1	239			
2	6518	1	239			
2	6519	1	239			
2	6520	1	239			
2	6521	1	239			
2	6522	1	239			
2	6523	1	239			
2	6524	1	239			
2	6525	1	239			
2	6526	1	239			
2	6527	1	239			
2	6528	1	239			
2	6529	1	256			
2	6530	1	256			
2	6531	1	256			
2	6532	1	256			
2	6533	1	256			
2	6534	1	256			
2	6535	1	256			
2	6536	1	256			
2	6537	1	256			
2	6538	1	256			
2	6539	1	256			
2	6540	1	256			
2	6541	1	256			
2	6542	1	256			
2	6543	1	256			
2	6544	1	256			
2	6545	1	273			
2	6546	1	273			
2	6547	1	273			
2	6548	1	273			
2	6549	1	273			
2	6550	1	273			
2	6551	1	273			
2	6552	1	273			
2	6553	1	273			
2	6554	1	273			
2	6555	1	273			
2	6556	1	273			
2	6557	1	273			
2	6558	1	273			
2	6559	1	273			
2	6560	1	273			
2	6561	1	290			
2	6562	1	290			
2	6563	1	290			
2	6564	1	290			
2	6565	1	290			
2	6566	1	290			
2	6567	1	290			
2	6568	1	290			
2	6569	1	290			
2	6570	1	290			
2	6571	1	290			
2	6572	1	290			
2	6573	1	290			
2	6574	1	290			
2	6575	1	290			
2	6576	1	290			
2	6577	1	307			
2	6578	1	307			
2	6579	1	307			
2	6580	1	307			
2	6581	1	307			
2	6582	1	307			
2	6583	1	307			
2	6584	1	307			
2	6585	1	307			
2	6586	1	307			
2	6587	1	307			
2	6588	1	307			
2	6589	1	307			
2	6590	1	307			
2	6591	1	307			
2	6592	1	307			
2	6593	1	324			
2	6594	1	324			
2	6595	1	324			
2	6596	1	324			
2	6597	1	324			
2	6598	1	324			
2	6599	1	324			
2	6600	1	324			
2	6601	1	324			
2	6602	1	324			
2	6603	1	324			
2	6604	1	324			
2	6605	1	324			
2	6606	1	324			
2	6607	1	324			
2	6608	1	324			
2	6609	1	341			
2	6610	1	341			
2	6611	1	341			
2	6612	1	341			
2	6613	1	341			
2	6614	1	341			
2	6615	1	341			
2	6616	1	341			
2	6617	1	341			
2	6618	1	341			
2	6619	1	341			
2	6620	1	341			
2	6621	1	341			
2	6622	1	341			
2	6623	1	341			
2	6624	1	341			
2	6625	1	358			
2	6626	1	358			
2	6627	1	358			
2	6628	1	358			
2	6629	1	358			
2	6630	1	358			
2	6631	1	358			
2	6632	1	358			
2	6633	1	358			
2	6634	1	358			
2	6635	1	358			
2	6636	1	358			
2	6637	1	358			
2	6638	1	358			
2	6639	1	358			
2	6640	1	358			
2	6641	1	375			
2	6642	1	375			
2	6643	1	375			
2	6644	1	375			
2	6645	1	375			
2	6646	1	375			
2	6647	1	375			
2	6648	1	375			
2	6649	1	375			
2	6650	1	375			
2	6651	1	375			
2	6652	1	375			
2	6653	1	375			
2	6654	1	375			
2	6655	1	375			
2	6656	1	375			
2	6657	1	392			
2	6658	1	392			
2	6659	1	392			
2	6660	1	392			
2	6661	1	392			
2	6662	1	392			
2	6663	1	392			
2	6664	1	392			
2	6665	1	392			
2	6666	1	392			
2	6667	1	392			
2	6668	1	392			
2	6669	1	392			
2	6670	1	392			
2	6671	1	392			
2	6672	1	392			
2	6673	1	409			
2	6674	1	409			
2	6675	1	409			
2	6676	1	409			
2	6677	1	409			
2	6678	1	409			
2	6679	1	409			
2	6680	1	409			
2	6681	1	409			
2	6682	1	409			
2	6683	1	409			
2	6684	1	409			
2	6685	1	409			
2	6686	1	409			
2	6687	1	409			
2	6688	1	409			
2	6689	1	426			
2	6690	1	426			
2	6691	1	426			
2	6692	1	426			
2	6693	1	426			
2	6694	1	426			
2	6695	1	426			
2	6696	1	426			
2	6697	1	426			
2	6698	1	426			
2	6699	1	426			
2	6700	1	426			
2	6701	1	426			
2	6702	1	426			
2	6703	1	426			
2	6704	1	426			
2	6705	1	443			
2	6706	1	443			
2	6707	1	443			
2	6708	1	443			
2	6709	1	443			
2	6710	1	443			
2	6711	1	443			
2	6712	1	443			
2	6713	1	443			
2	6714	1	443			
2	6715	1	443			
2	6716	1	443			
2	6717	1	443			
2	6718	1	443			
2	6719	1	443			
2	6720	1	443			
2	6721	1	460			
2	6722	1	460			
2	6723	1	460			
2	6724	1	460			
2	6725	1	460			
2	6726	1	460			
2	6727	1	460			
2	6728	1	460			
2	6729	1	460			
2	6730	1	460			
2	6731	1	460			
2	6732	1	460			
2	6733	1	460			
2	6734	1	460			
2	6735	1	460			
2	6736	1	460			
2	6737	1	477			
2	6738	1	477			
2	6739	1	477			
2	6740	1	477			
2	6741	1	477			
2	6742	1	477			
2	6743	1	477			
2	6744	1	477			
2	6745	1	477			
2	6746	1	477			
2	6747	1	477			
2	6748	1	477			
2	6749	1	477			
2	6750	1	477			
2	6751	1	477			
2	6752	1	477			
2	6753	1	494			
2	6754	1	494			
2	6755	1	494			
2	6756	1	494			
2	6757	1	494			
2	6758	1	494			
2	6759	1	494			
2	6760	1	494			
2	6761	1	494			
2	6762	1	494			
2	6763	1	494			
2	6764	1	494			
2	6765	1	494			
2	6766	1	494			
2	6767	1	494			
2	6768	1	494			
2	6769	1	511			
2	6770	1	511			
2	6771	1	511			
2	6772	1	511			
2	6773	1	511			
2	6774	1	511			
2	6775	1	511			
2	6776	1	511			
2	6777	1	511			
2	6778	1	511			
2	6779	1	511			
2	6780	1	511			
2	6781	1	511			
2	6782	1	511			
2	6783	1	511			
2	6784	1	511			
2	6785	1	528			
2	6786	1	528			
2	6787	1	528			
2	6788	1	528			
2	6789	1	528			
2	6790	1	528			
2	6791	1	528			
2	6792	1	528			
2	6793	1	528			
2	6794	1	528			
2	6795	1	528			
2	6796	1	528			
2	6797	1	528			
2	6798	1	528			
2	6799	1	528			
2	6800	1	528			
2	6801	1	546			
2	6802	1	546			
2	6803	1	549			
2	6804	1	549			
2	6805	1	552			
2	6806	1	552			
2	6807	1	555			
2	6808	1	555			
2	6809	1	558			
2	6810	1	558			
2	6811	1	561			
2	6812	1	561			
2	6813	1	564			
2	6814	1	564			
2	6815	1	567			
2	6816	1	567			
2	6817	1	570			
2	6818	1	570			
2	6819	1	573			
2	6820	1	573			
2	6821	1	576			
2	6822	1	576			
2	6823	1	579			
2	6824	1	579			
2	6825	1	582			
2	6826	1	582			
2	6827	1	585			
2	6828	1	585			
2	6829	1	588			
2	6830	1	588			
2	6831	1	591			
2	6832	1	591			
2	6833	1	594			
2	6834	1	594			
2	6835	1	597			
2	6836	1	597			
2	6837	1	600			
2	6838	1	600			
2	6839	1	603			
2	6840	1	603			
2	6841	1	606			
2	6842	1	606			
2	6843	1	609			
2	6844	1	609			
2	6845	1	612			
2	6846	1	612			
2	6847	1	615			
2	6848	1	615			
2	6849	1	618			
2	6850	1	618			
2	6851	1	621			
2	6852	1	621			
2	6853	1	624			
2	6854	1	624			
2	6855	1	627			
2	6856	1	627			
2	6857	1	630			
2	6858	1	630			
2	6859	1	633			
2	6860	1	633			
2	6861	1	636			
2	6862	1	636			
2	6863	1	639			
2	6864	1	639			
2	6865	1	642			
2	6866	1	642			
2	6867	1	645			
2	6868	1	645			
2	6869	1	648			
2	6870	1	648			
2	6871	1	651			
2	6872	1	651			
2	6873	1	654			
2	6874	1	654			
2	6875	1	657			
2	6876	1	657			
2	6877	1	660			
2	6878	1	660			
2	6879	1	663			
2	6880	1	663			
2	6881	1	666			
2	6882	1	666			
2	6883	1	669			
2	6884	1	669			
2	6885	1	672			
2	6886	1	672			
2	6887	1	675			
2	6888	1	675			
2	6889	1	678			
2	6890	1	678			
2	6891	1	681			
2	6892	1	681			
2	6893	1	684			
2	6894	1	684			
2	6895	1	687			
2	6896	1	687			
2	6897	1	690			
2	6898	1	690			
2	6899	1	693			
2	6900	1	693			
2	6901	1	696			
2	6902	1	696			
2	6903	1	699			
2	6904	1	699			
2	6905	1	702			
2	6906	1	702			
2	6907	1	705			
2	6908	1	705			
2	6909	1	708			
2	6910	1	708			
2	6911	1	711			
2	6912	1	711			
2	6913	1	714			
2	6914	1	714			
2	6915	1	717			
2	6916	1	717			
2	6917	1	720			
2	6918	1	720			
2	6919	1	723			
2	6920	1	723			
2	6921	1	726			
2	6922	1	726			
2	6923	1	729			
2	6924	1	729			
2	6925	1	732			
2	6926	1	732			
2	6927	1	735			
2	6928	1	735			
2	6929	1	738			
2	6930	1	738			
2	6931	1	741			
2	6932	1	741			
2	6933	1	744			
2	6934	1	744			
2	6935	1	747			
2	6936	1	747			
2	6937	1	750			
2	6938	1	750			
2	6939	1	753			
2	6940	1	753			
2	6941	1	756			
2	6942	1	756			
2	6943	1	759			
2	6944	1	759			
2	6945	1	762			
2	6946	1	762			
2	6947	1	765			
2	6948	1	765			
2	6949	1	768			
2	6950	1	768			
2	6951	1	771			
2	6952	1	771			
2	6953	1	774			
2	6954	1	774			
2	6955	1	777			
2	6956	1	777			
2	6957	1	780			
2	6958	1	780			
2	6959	1	783			
2	6960	1	783			
2	6961	1	786			
2	6962	1	786			
2	6963	1	789			
2	6964	1	789			
2	6965	1	792			
2	6966	1	792			
2	6967	1	795			
2	6968	1	795			
2	6969	1	798			
2	6970	1	798			
2	6971	1	801			
2	6972	1	801			
2	6973	1	804			
2	6974	1	804			
2	6975	1	807			
2	6976	1	807			
2	6977	1	810			
2	6978	1	810			
2	6979	1	813			
2	6980	1	813			
2	6981	1	816			
2	6982	1	816			
2	6983	1	819			
2	6984	1	819			
2	6985	1	822			
2	6986	1	822			
2	6987	1	825			
2	6988	1	825			
2	6989	1	828			
2	6990	1	828			
2	6991	1	831			
2	6992	1	831			
2	6993	1	834			
2	6994	1	834			
2	6995	1	837			
2	6996	1	837			
2	6997	1	840			
2	6998	1	840			
2	6999	1	843			
2	7000	1	843			
2	7001	1	846			
2	7002	1	846			
2	7003	1	849			
2	7004	1	849			
2	7005	1	852			
2	7006	1	852			
2	7007	1	855			
2	7008	1	855			
2	7009	1	858			
2	7010	1	858			
2	7011	1	861			
2	7012	1	861			
2	7013	1	864			
2	7014	1	864			
2	7015	1	867			
2	7016	1	867			
2	7017	1	870			
2	7018	1	870			
2	7019	1	873			
2	7020	1	873			
2	7021	1	876			
2	7022	1	876			
2	7023	1	879			
2	7024	1	879			
2	7025	1	882			
2	7026	1	882			
2	7027	1	885			
2	7028	1	885			
2	7029	1	888			
2	7030	1	888			
2	7031	1	891			
2	7032	1	891			
2	7033	1	894			
2	7034	1	894			
2	7035	1	897			
2	7036	1	897			
2	7037	1	900			
2	7038	1	900			
2	7039	1	903			
2	7040	1	903			
2	7041	1	906			
2	7042	1	906			
2	7043	1	909			
2	7044	1	909			
2	7045	1	912			
2	7046	1	912			
2	7047	1	915			
2	7048	1	915			
2	7049	1	918			
2	7050	1	918			
2	7051	1	921			
2	7052	1	921			
2	7053	1	924			
2	7054	1	924			
2	7055	1	927			
2	7056	1	927			
2	7057	1	930			
2	7058	1	930			
2	7059	1	933			
2	7060	1	933			
2	7061	1	936			
2	7062	1	936			
2	7063	1	939			
2	7064	1	939			
2	7065	1	942			
2	7066	1	942			
2	7067	1	945			
2	7068	1	945			
2	7069	1	948			
2	7070	1	948			
2	7071	1	951			
2	7072	1	951			
2	7073	1	954			
2	7074	1	954			
2	7075	1	957			
2	7076	1	957			
2	7077	1	960			
2	7078	1	960			
2	7079	1	963			
2	7080	1	963			
2	7081	1	966			
2	7082	1	966			
2	7083	1	969			
2	7084	1	969			
2	7085	1	972			
2	7086	1	972			
2	7087	1	975			
2	7088	1	975			
2	7089	1	978			
2	7090	1	978			
2	7091	1	981			
2	7092	1	981			
2	7093	1	984			
2	7094	1	984			
2	7095	1	987			
2	7096	1	987			
2	7097	1	990			
2	7098	1	990			
2	7099	1	993			
2	7100	1	993			
2	7101	1	996			
2	7102	1	996			
2	7103	1	999			
2	7104	1	999			
2	7105	1	1002			
2	7106	1	1002			
2	7107	1	1005			
2	7108	1	1005			
2	7109	1	1008			
2	7110	1	1008			
2	7111	1	1011			
2	7112	1	1011			
2	7113	1	1014			
2	7114	1	1014			
2	7115	1	1017			
2	7116	1	1017			
2	7117	1	1020			
2	7118	1	1020			
2	7119	1	1023			
2	7120	1	1023			
2	7121	1	1026			
2	7122	1	1026			
2	7123	1	1029			
2	7124	1	1029			
2	7125	1	1032			
2	7126	1	1032			
2	7127	1	1035			
2	7128	1	1035			
2	7129	1	1038			
2	7130	1	1038			
2	7131	1	1041			
2	7132	1	1041			
2	7133	1	1044			
2	7134	1	1044			
2	7135	1	1047			
2	7136	1	1047			
2	7137	1	1050			
2	7138	1	1050			
2	7139	1	1053			
2	7140	1	1053			
2	7141	1	1056			
2	7142	1	1056			
2	7143	1	1059			
2	7144	1	1059			
2	7145	1	1062			
2	7146	1	1062			
2	7147	1	1065			
2	7148	1	1065			
2	7149	1	1068			
2	7150	1	1068			
2	7151	1	1071			
2	7152	1	1071			
2	7153	1	1074			
2	7154	1	1074			
2	7155	1	1077			
2	7156	1	1077			
2	7157	1	1080			
2	7158	1	1080			
2	7159	1	1083			
2	7160	1	1083			
2	7161	1	1086			
2	7162	1	1086			
2	7163	1	1089			
2	7164	1	1089			
2	7165	1	1092			
2	7166	1	1092			
2	7167	1	1095			
2	7168	1	1095			
2	7169	1	1098			
2	7170	1	1098			
2	7171	1	1101			
2	7172	1	1101			
2	7173	1	1104			
2	7174	1	1104			
2	7175	1	1107			
2	7176	1	1107			
2	7177	1	1110			
2	7178	1	1110			
2	7179	1	1113			
2	7180	1	1113			
2	7181	1	1116			
2	7182	1	1116			
2	7183	1	1119			
2	7184	1	1119			
2	7185	1	1122			
2	7186	1	1122			
2	7187	1	1125			
2	7188	1	1125			
2	7189	1	1128			
2	7190	1	1128			
2	7191	1	1131			
2	7192	1	1131			
2	7193	1	1134			
2	7194	1	1134			
2	7195	1	1137			
2	7196	1	1137			
2	7197	1	1140			
2	7198	1	1140			
2	7199	1	1143			
2	7200	1	1143			
2	7201	1	1146			
2	7202	1	1146			
2	7203	1	1149			
2	7204	1	1149			
2	7205	1	1152			
2	7206	1	1152			
2	7207	1	1155			
2	7208	1	1155			
2	7209	1	1158			
2	7210	1	1158			
2	7211	1	1161			
2	7212	1	1161			
2	7213	1	1164			
2	7214	1	1164			
2	7215	1	1167			
2	7216	1	1167			
2	7217	1	1170			
2	7218	1	1170			
2	7219	1	1173			
2	7220	1	1173			
2	7221	1	1176			
2	7222	1	1176			
2	7223	1	1179			
2	7224	1	1179			
2	7225	1	1182			
2	7226	1	1182			
2	7227	1	1185			
2	7228	1	1185			
2	7229	1	1188			
2	7230	1	1188			
2	7231	1	1191			
2	7232	1	1191			
2	7233	1	1194			
2	7234	1	1194			
2	7235	1	1197			
2	7236	1	1197			
2	7237	1	1200			
2	7238	1	1200			
2	7239	1	1203			
2	7240	1	1203			
2	7241	1	1206			
2	7242	1	1206			
2	7243	1	1209			
2	7244	1	1209			
2	7245	1	1212			
2	7246	1	1212			
2	7247	1	1215			
2	7248	1	1215			
2	7249	1	1218			
2	7250	1	1218			
2	7251	1	1221			
2	7252	1	1221			
2	7253	1	1224			
2	7254	1	1224			
2	7255	1	1227			
2	7256	1	1227			
2	7257	1	1230			
2	7258	1	1230			
2	7259	1	1233			
2	7260	1	1233			
2	7261	1	1236			
2	7262	1	1236			
2	7263	1	1239			
2	7264	1	1239			
2	7265	1	1242			
2	7266	1	1242			
2	7267	1	1245			
2	7268	1	1245			
2	7269	1	1248			
2	7270	1	1248			
2	7271	1	1251			
2	7272	1	1251			
2	7273	1	1254			
2	7274	1	1254			
2	7275	1	1257			
2	7276	1	1257			
2	7277	1	1260			
2	7278	1	1260			
2	7279	1	1263			
2	7280	1	1263			
2	7281	1	1266			
2	7282	1	1266			
2	7283	1	1269			
2	7284	1	1269			
2	7285	1	1272			
2	7286	1	1272			
2	7287	1	1275			
2	7288	1	1275			
2	7289	1	1278			
2	7290	1	1278			
2	7291	1	1281			
2	7292	1	1281			
2	7293	1	1284			
2	7294	1	1284			
2	7295	1	1287			
2	7296	1	1287			
2	7297	1	1290			
2	7298	1	1290			
2	7299	1	1293			
2	7300	1	1293			
2	7301	1	1296			
2	7302	1	1296			
2	7303	1	1299			
2	7304	1	1299			
2	7305	1	1302			
2	7306	1	1302			
2	7307	1	1305			
2	7308	1	1305			
2	7309	1	1308			
2	7310	1	1308			
2	7311	1	1311			
2	7312	1	1311			
2	7313	1	1311			
2	7314	1	1315			
2	7315	1	1315			
2	7316	1	1315			
2	7317	1	1319			
2	7318	1	1319			
2	7319	1	1319			
2	7320	1	1323			
2	7321	1	1323			
2	7322	1	1323			
2	7323	1	1327			
2	7324	1	1327			
2	7325	1	1327			
2	7326	1	1331			
2	7327	1	1331			
2	7328	1	1331			
2	7329	1	1335			
2	7330	1	1335			
2	7331	1	1335			
2	7332	1	1339			
2	7333	1	1339			
2	7334	1	1339			
2	7335	1	1343			
2	7336	1	1343			
2	7337	1	1343			
2	7338	1	1347			
2	7339	1	1347			
2	7340	1	1347			
2	7341	1	1351			
2	7342	1	1351			
2	7343	1	1351			
2	7344	1	1355			
2	7345	1	1355			
2	7346	1	1355			
2	7347	1	1359			
2	7348	1	1359			
2	7349	1	1359			
2	7350	1	1363			
2	7351	1	1363			
2	7352	1	1363			
2	7353	1	1367			
2	7354	1	1367			
2	7355	1	1367			
2	7356	1	1401			
2	7357	1	1401			
2	7358	1	1404			
2	7359	1	1404			
2	7360	1	1407			
2	7361	1	1407			
2	7362	1	1410			
2	7363	1	1410			
2	7364	1	1413			
2	7365	1	1413			
2	7366	1	1416			
2	7367	1	1416			
2	7368	1	1419			
2	7369	1	1419			
2	7370	1	1422			
2	7371	1	1422			
2	7372	1	1425			
2	7373	1	1425			
2	7374	1	1428			
2	7375	1	1428			
2	7376	1	1431			
2	7377	1	1431			
2	7378	1	1434			
2	7379	1	1434			
2	7380	1	1437			
2	7381	1	1437			
2	7382	1	1440			
2	7383	1	1440			
2	7384	1	1443			
2	7385	1	1443			
2	7386	1	1446			
2	7387	1	1446			
2	7388	1	1446			
2	7389	1	1450			
2	7390	1	1450			
2	7391	1	1450			
2	7392	1	1454			
2	7393	1	1454			
2	7394	1	1454			
2	7395	1	1458			
2	7396	1	1458			
2	7397	1	1458			
2	7398	1	1462			
2	7399	1	1462			
2	7400	1	1462			
2	7401	1	1466			
2	7402	1	1466			
2	7403	1	1466			
2	7404	1	1470			
2	7405	1	1470			
2	7406	1	1470			
2	7407	1	1474			
2	7408	1	1474			
2	7409	1	1474			
2	7410	1	1478			
2	7411	1	1478			
2	7412	1	1478			
2	7413	1	1482			
2	7414	1	1482			
2	7415	1	1482			
2	7416	1	1486			
2	7417	1	1486			
2	7418	1	1486			
2	7419	1	1490			
2	7420	1	1490			
2	7421	1	1490			
2	7422	1	1494			
2	7423	1	1494			
2	7424	1	1494			
2	7425	1	1498			
2	7426	1	1498			
2	7427	1	1498			
2	7428	1	1502			
2	7429	1	1502			
2	7430	1	1502			
2	7431	1	1508			
2	7432	1	1508			
2	7433	1	1513			
2	7434	1	1513			
2	7435	1	1518			
2	7436	1	1518			
2	7437	1	1523			
2	7438	1	1523			
2	7439	1	1528			
2	7440	1	1528			
2	7441	1	1533			
2	7442	1	1533			
2	7443	1	1538			
2	7444	1	1538			
2	7445	1	1543			
2	7446	1	1543			
2	7447	1	1548			
2	7448	1	1548			
2	7449	1	1553			
2	7450	1	1553			
2	7451	1	1558			
2	7452	1	1558			
2	7453	1	1563			
2	7454	1	1563			
2	7455	1	1568			
2	7456	1	1568			
2	7457	1	1573			
2	7458	1	1573			
2	7459	1	1578			
2	7460	1	1578			
2	7461	1	1582			
2	7462	1	1582			
2	7463	1	1585			
2	7464	1	1585			
2	7465	1	1588			
2	7466	1	1588			
2	7467	1	1591			
2	7468	1	1591			
2	7469	1	1594			
2	7470	1	1594			
2	7471	1	1597			
2	7472	1	1597			
2	7473	1	1600			
2	7474	1	1600			
2	7475	1	1603			
2	7476	1	1603			
2	7477	1	1606			
2	7478	1	1606			
2	7479	1	1609			
2	7480	1	1609			
2	7481	1	1612			
2	7482	1	1612			
2	7483	1	1615			
2	7484	1	1615			
2	7485	1	1618			
2	7486	1	1618			
2	7487	1	1621			
2	7488	1	1621			
2	7489	1	1624			
2	7490	1	1624			
2	7491	1	1624			
2	7492	1	1628			
2	7493	1	1628			
2	7494	1	1628			
2	7495	1	1632			
2	7496	1	1632			
2	7497	1	1632			
2	7498	1	1636			
2	7499	1	1636			
2	7500	1	1636			
2	7501	1	1640			
2	7502	1	1640			
2	7503	1	1640			
2	7504	1	1644			
2	7505	1	1644			
2	7506	1	1644			
2	7507	1	1648			
2	7508	1	1648			
2	7509	1	1648			
2	7510	1	1652			
2	7511	1	1652			
2	7512	1	1652			
2	7513	1	1656			
2	7514	1	1656			
2	7515	1	1656			
2	7516	1	1660			
2	7517	1	1660			
2	7518	1	1660			
2	7519	1	1664			
2	7520	1	1664			
2	7521	1	1664			
2	7522	1	1668			
2	7523	1	1668			
2	7524	1	1668			
2	7525	1	1672			
2	7526	1	1672			
2	7527	1	1672			
2	7528	1	1676			
2	7529	1	1676			
2	7530	1	1676			
2	7531	1	1680			
2	7532	1	1680			
2	7533	1	1680			
2	7534	1	1714			
2	7535	1	1714			
2	7536	1	1717			
2	7537	1	1717			
2	7538	1	1720			
2	7539	1	1720			
2	7540	1	1723			
2	7541	1	1723			
2	7542	1	1726			
2	7543	1	1726			
2	7544	1	1729			
2	7545	1	1729			
2	7546	1	1732			
2	7547	1	1732			
2	7548	1	1735			
2	7549	1	1735			
2	7550	1	1738			
2	7551	1	1738			
2	7552	1	1741			
2	7553	1	1741			
2	7554	1	1744			
2	7555	1	1744			
2	7556	1	1747			
2	7557	1	1747			
2	7558	1	1750			
2	7559	1	1750			
2	7560	1	1753			
2	7561	1	1753			
2	7562	1	1756			
2	7563	1	1756			
2	7564	1	1759			
2	7565	1	1759			
2	7566	1	1759			
2	7567	1	1763			
2	7568	1	1763			
2	7569	1	1763			
2	7570	1	1767			
2	7571	1	1767			
2	7572	1	1767			
2	7573	1	1771			
2	7574	1	1771			
2	7575	1	1771			
2	7576	1	1775			
2	7577	1	1775			
2	7578	1	1775			
2	7579	1	1779			
2	7580	1	1779			
2	7581	1	1779			
2	7582	1	1783			
2	7583	1	1783			
2	7584	1	1783			
2	7585	1	1787			
2	7586	1	1787			
2	7587	1	1787			
2	7588	1	1791			
2	7589	1	1791			
2	7590	1	1791			
2	7591	1	1795			
2	7592	1	1795			
2	7593	1	1795			
2	7594	1	1799			
2	7595	1	1799			
2	7596	1	1799			
2	7597	1	1803			
2	7598	1	1803			
2	7599	1	1803			
2	7600	1	1807			
2	7601	1	1807			
2	7602	1	1807			
2	7603	1	1811			
2	7604	1	1811			
2	7605	1	1811			
2	7606	1	1815			
2	7607	1	1815			
2	7608	1	1815			
2	7609	1	1821			
2	7610	1	1821			
2	7611	1	1826			
2	7612	1	1826			
2	7613	1	1831			
2	7614	1	1831			
2	7615	1	1836			
2	7616	1	1836			
2	7617	1	1841			
2	7618	1	1841			
2	7619	1	1846			
2	7620	1	1846			
2	7621	1	1851			
2	7622	1	1851			
2	7623	1	1856			
2	7624	1	1856			
2	7625	1	1861			
2	7626	1	1861			
2	7627	1	1866			
2	7628	1	1866			
2	7629	1	1871			
2	7630	1	1871			
2	7631	1	1876			
2	7632	1	1876			
2	7633	1	1881			
2	7634	1	1881			
2	7635	1	1886			
2	7636	1	1886			
2	7637	1	1891			
2	7638	1	1891			
2	7639	1	1894			
2	7640	1	1894			
2	7641	1	1897			
2	7642	1	1897			
2	7643	1	1897			
2	7644	1	1902			
2	7645	1	1902			
2	7646	1	1905			
2	7647	1	1905			
2	7648	1	1908			
2	7649	1	1908			
2	7650	1	1911			
2	7651	1	1911			
2	7652	1	1914			
2	7653	1	1914			
2	7654	1	1917			
2	7655	1	1917			
2	7656	1	1920			
2	7657	1	1920			
2	7658	1	1923			
2	7659	1	1923			
2	7660	1	1926			
2	7661	1	1926			
2	7662	1	1929			
2	7663	1	1929			
2	7664	1	1932			
2	7665	1	1932			
2	7666	1	1935			
2	7667	1	1935			
2	7668	1	1938			
2	7669	1	1938			
2	7670	1	1941			
2	7671	1	1941			
2	7672	1	1941			
2	7673	1	1947			
2	7674	1	1947			
2	7675	1	1947			
2	7676	1	1951			
2	7677	1	1951			
2	7678	1	1951			
2	7679	1	1955			
2	7680	1	1955			
2	7681	1	1955			
2	7682	1	1959			
2	7683	1	1959			
2	7684	1	1959			
2	7685	1	1963			
2	7686	1	1963			
2	7687	1	1963			
2	7688	1	1967			
2	7689	1	1967			
2	7690	1	1967			
2	7691	1	1971			
2	7692	1	1971			
2	7693	1	1971			
2	7694	1	1975			
2	7695	1	1975			
2	7696	1	1975			
2	7697	1	1979			
2	7698	1	1979			
2	7699	1	1979			
2	7700	1	1983			
2	7701	1	1983			
2	7702	1	1983			
2	7703	1	1987			
2	7704	1	1987			
2	7705	1	1987			
2	7706	1	1991			
2	7707	1	1991			
2	7708	1	1991			
2	7709	1	1995			
2	7710	1	1995			
2	7711	1	1995			
2	7712	1	2001			
2	7713	1	2001			
2	7714	1	2030			
2	7715	1	2030			
2	7716	1	2033			
2	7717	1	2033			
2	7718	1	2033			
2	7719	1	2037			
2	7720	1	2037			
2	7721	1	2040			
2	7722	1	2040			
2	7723	1	2043			
2	7724	1	2043			
2	7725	1	2046			
2	7726	1	2046			
2	7727	1	2049			
2	7728	1	2049			
2	7729	1	2052			
2	7730	1	2052			
2	7731	1	2055			
2	7732	1	2055			
2	7733	1	2058			
2	7734	1	2058			
2	7735	1	2061			
2	7736	1	2061			
2	7737	1	2064			
2	7738	1	2064			
2	7739	1	2067			
2	7740	1	2067			
2	7741	1	2070			
2	7742	1	2070			
2	7743	1	2073			
2	7744	1	2073			
2	7745	1	2076			
2	7746	1	2076			
2	7747	1	2076			
2	7748	1	2082			
2	7749	1	2082			
2	7750	1	2085			
2	7751	1	2085			
2	7752	1	2085			
2	7753	1	2089			
2	7754	1	2089			
2	7755	1	2089			
2	7756	1	2093			
2	7757	1	2093			
2	7758	1	2093			
2	7759	1	2097			
2	7760	1	2097			
2	7761	1	2097			
2	7762	1	2101			
2	7763	1	2101			
2	7764	1	2101			
2	7765	1	2105			
2	7766	1	2105			
2	7767	1	2105			
2	7768	1	2109			
2	7769	1	2109			
2	7770	1	2109			
2	7771	1	2113			
2	7772	1	2113			
2	7773	1	2113			
2	7774	1	2117			
2	7775	1	2117			
2	7776	1	2117			
2	7777	1	2121			
2	7778	1	2121			
2	7779	1	2121			
2	7780	1	2125			
2	7781	1	2125			
2	7782	1	2125			
2	7783	1	2129			
2	7784	1	2129			
2	7785	1	2129			
2	7786	1	2133			
2	7787	1	2133			
2	7788	1	2133			
2	7789	1	2139			
2	7790	1	2139			
2	7791	1	2142			
2	7792	1	2142			
2	7793	1	2145			
2	7794	1	2145			
2	7795	1	2145			
2	7796	1	2151			
2	7797	1	2151			
2	7798	1	2156			
2	7799	1	2156			
2	7800	1	2161			
2	7801	1	2161			
2	7802	1	2166			
2	7803	1	2166			
2	7804	1	2171			
2	7805	1	2171			
2	7806	1	2176			
2	7807	1	2176			
2	7808	1	2181			
2	7809	1	2181			
2	7810	1	2186			
2	7811	1	2186			
2	7812	1	2191			
2	7813	1	2191			
2	7814	1	2196			
2	7815	1	2196			
2	7816	1	2201			
2	7817	1	2201			
2	7818	1	2206			
2	7819	1	2206			
2	7820	1	2211			
2	7821	1	2211			
2	7822	1	2214			
2	7823	1	2214			
2	7824	1	2217			
2	7825	1	2217			
2	7826	1	2217			
2	7827	1	2224			
2	7828	1	2224			
2	7829	1	2227			
2	7830	1	2227			
2	7831	1	2230			
2	7832	1	2230			
2	7833	1	2233			
2	7834	1	2233			
2	7835	1	2236			
2	7836	1	2236			
2	7837	1	2239			
2	7838	1	2239			
2	7839	1	2242			
2	7840	1	2242			
2	7841	1	2245			
2	7842	1	2245			
2	7843	1	2248			
2	7844	1	2248			
2	7845	1	2251			
2	7846	1	2251			
2	7847	1	2254			
2	7848	1	2254			
2	7849	1	2257			
2	7850	1	2257			
2	7851	1	2260			
2	7852	1	2260			
2	7853	1	2260			
2	7854	1	2266			
2	7855	1	2266			
2	7856	1	2269			
2	7857	1	2269			
2	7858	1	2269			
2	7859	1	2273			
2	7860	1	2273			
2	7861	1	2273			
2	7862	1	2277			
2	7863	1	2277			
2	7864	1	2277			
2	7865	1	2281			
2	7866	1	2281			
2	7867	1	2281			
2	7868	1	2285			
2	7869	1	2285			
2	7870	1	2285			
2	7871	1	2289			
2	7872	1	2289			
2	7873	1	2289			
2	7874	1	2293			
2	7875	1	2293			
2	7876	1	2293			
2	7877	1	2297			
2	7878	1	2297			
2	7879	1	2297			
2	7880	1	2301			
2	7881	1	2301			
2	7882	1	2301			
2	7883	1	2305			
2	7884	1	2305			
2	7885	1	2305			
2	7886	1	2309			
2	7887	1	2309			
2	7888	1	2309			
2	7889	1	2313			
2	7890	1	2313			
2	7891	1	2313			
2	7892	1	2319			
2	7893	1	2319			
2	7894	1	2322			
2	7895	1	2322			
2	7896	1	2322			
2	7897	1	2350			
2	7898	1	2350			
2	7899	1	2353			
2	7900	1	2353			
2	7901	1	2353			
2	7902	1	2359			
2	7903	1	2359			
2	7904	1	2362			
2	7905	1	2362			
2	7906	1	2365			
2	7907	1	2365			
2	7908	1	2368			
2	7909	1	2368			
2	7910	1	2371			
2	7911	1	2371			
2	7912	1	2374			
2	7913	1	2374			
2	7914	1	2377			
2	7915	1	2377			
2	7916	1	2380			
2	7917	1	2380			
2	7918	1	2383			
2	7919	1	2383			
2	7920	1	2386			
2	7921	1	2386			
2	7922	1	2389			
2	7923	1	2389			
2	7924	1	2392			
2	7925	1	2392			
2	7926	1	2395			
2	7927	1	2395			
2	7928	1	2398			
2	7929	1	2398			
2	7930	1	2398			
2	7931	1	2404			
2	7932	1	2404			
2	7933	1	2407			
2	7934	1	2407			
2	7935	1	2410			
2	7936	1	2410			
2	7937	1	2410			
2	7938	1	2414			
2	7939	1	2414			
2	7940	1	2414			
2	7941	1	2418			
2	7942	1	2418			
2	7943	1	2418			
2	7944	1	2422			
2	7945	1	2422			
2	7946	1	2422			
2	7947	1	2426			
2	7948	1	2426			
2	7949	1	2426			
2	7950	1	2430			
2	7951	1	2430			
2	7952	1	2430			
2	7953	1	2434			
2	7954	1	2434			
2	7955	1	2434			
2	7956	1	2438			
2	7957	1	2438			
2	7958	1	2438			
2	7959	1	2442			
2	7960	1	2442			
2	7961	1	2442			
2	7962	1	2446			
2	7963	1	2446			
2	7964	1	2446			
2	7965	1	2450			
2	7966	1	2450			
2	7967	1	2450			
2	7968	1	2454			
2	7969	1	2454			
2	7970	1	2454			
2	7971	1	2458			
2	7972	1	2458			
2	7973	1	2458			
2	7974	1	2464			
2	7975	1	2464			
2	7976	1	2467			
2	7977	1	2467			
2	7978	1	2470			
2	7979	1	2470			
2	7980	1	2470			
2	7981	1	2478			
2	7982	1	2478			
2	7983	1	2483			
2	7984	1	2483			
2	7985	1	2488			
2	7986	1	2488			
2	7987	1	2493			
2	7988	1	2493			
2	7989	1	2498			
2	7990	1	2498			
2	7991	1	2503			
2	7992	1	2503			
2	7993	1	2508			
2	7994	1	2508			
2	7995	1	2513			
2	7996	1	2513			
2	7997	1	2518			
2	7998	1	2518			
2	7999	1	2523			
2	8000	1	2523			
2	8001	1	2528			
2	8002	1	2528			
2	8003	1	2533			
2	8004	1	2533			
2	8005	1	2536			
2	8006	1	2536			
2	8007	1	2539			
2	8008	1	2539			
2	8009	1	2539			
2	8010	1	2545			
2	8011	1	2545			
2	8012	1	2549			
2	8013	1	2549			
2	8014	1	2552			
2	8015	1	2552			
2	8016	1	2555			
2	8017	1	2555			
2	8018	1	2558			
2	8019	1	2558			
2	8020	1	2561			
2	8021	1	2561			
2	8022	1	2564			
2	8023	1	2564			
2	8024	1	2567			
2	8025	1	2567			
2	8026	1	2570			
2	8027	1	2570			
2	8028	1	2573			
2	8029	1	2573			
2	8030	1	2576			
2	8031	1	2576			
2	8032	1	2579			
2	8033	1	2579			
2	8034	1	2582			
2	8035	1	2582			
2	8036	1	2582			
2	8037	1	2588			
2	8038	1	2588			
2	8039	1	2591			
2	8040	1	2591			
2	8041	1	2591			
2	8042	1	2595			
2	8043	1	2595			
2	8044	1	2595			
2	8045	1	2599			
2	8046	1	2599			
2	8047	1	2599			
2	8048	1	2603			
2	8049	1	2603			
2	8050	1	2603			
2	8051	1	2607			
2	8052	1	2607			
2	8053	1	2607			
2	8054	1	2611			
2	8055	1	2611			
2	8056	1	2611			
2	8057	1	2615			
2	8058	1	2615			
2	8059	1	2615			
2	8060	1	2619			
2	8061	1	2619			
2	8062	1	2619			
2	8063	1	2623			
2	8064	1	2623			
2	8065	1	2623			
2	8066	1	2627			
2	8067	1	2627			
2	8068	1	2627			
2	8069	1	2631			
2	8070	1	2631			
2	8071	1	2631			
2	8072	1	2635			
2	8073	1	2635			
2	8074	1	2635			
2	8075	1	2641			
2	8076	1	2641			
2	8077	1	2644			
2	8078	1	2644			
2	8079	1	2644			
2	8080	1	2650			
2	8081	1	2650			
2	8082	1	2675			
2	8083	1	2675			
2	8084	1	2678			
2	8085	1	2678			
2	8086	1	2678			
2	8087	1	2684			
2	8088	1	2684			
2	8089	1	2687			
2	8090	1	2687			
2	8091	1	2690			
2	8092	1	2690			
2	8093	1	2690			
2	8094	1	2694			
2	8095	1	2694			
2	8096	1	2697			
2	8097	1	2697			
2	8098	1	2700			
2	8099	1	2700			
2	8100	1	2703			
2	8101	1	2703			
2	8102	1	2706			
2	8103	1	2706			
2	8104	1	2709			
2	8105	1	2709			
2	8106	1	2712			
2	8107	1	2712			
2	8108	1	2715			
2	8109	1	2715			
2	8110	1	2718			
2	8111	1	2718			
2	8112	1	2721			
2	8113	1	2721			
2	8114	1	2724			
2	8115	1	2724			
2	8116	1	2727			
2	8117	1	2727			
2	8118	1	2727			
2	8119	1	2733			
2	8120	1	2733			
2	8121	1	2736			
2	8122	1	2736			
2	8123	1	2739			
2	8124	1	2739			
2	8125	1	2739			
2	8126	1	2745			
2	8127	1	2745			
2	8128	1	2745			
2	8129	1	2749			
2	8130	1	2749			
2	8131	1	2749			
2	8132	1	2753			
2	8133	1	2753			
2	8134	1	2753			
2	8135	1	2757			
2	8136	1	2757			
2	8137	1	2757			
2	8138	1	2761			
2	8139	1	2761			
2	8140	1	2761			
2	8141	1	2765			
2	8142	1	2765			
2	8143	1	2765			
2	8144	1	2769			
2	8145	1	2769			
2	8146	1	2769			
2	8147	1	2773			
2	8148	1	2773			
2	8149	1	2773			
2	8150	1	2777			
2	8151	1	2777			
2	8152	1	2777			
2	8153	1	2781			
2	8154	1	2781			
2	8155	1	2781			
2	8156	1	2785			
2	8157	1	2785			
2	8158	1	2785			
2	8159	1	2791			
2	8160	1	2791			
2	8161	1	2794			
2	8162	1	2794			
2	8163	1	2797			
2	8164	1	2797			
2	8165	1	2797			
2	8166	1	2803			
2	8167	1	2803			
2	8168	1	2808			
2	8169	1	2808			
2	8170	1	2813			
2	8171	1	2813			
2	8172	1	2818			
2	8173	1	2818			
2	8174	1	2823			
2	8175	1	2823			
2	8176	1	2828			
2	8177	1	2828			
2	8178	1	2833			
2	8179	1	2833			
2	8180	1	2838			
2	8181	1	2838			
2	8182	1	2843			
2	8183	1	2843			
2	8184	1	2848			
2	8185	1	2848			
2	8186	1	2853			
2	8187	1	2853			
2	8188	1	2858			
2	8189	1	2858			
2	8190	1	2861			
2	8191	1	2861			
2	8192	1	2864			
2	8193	1	2864			
2	8194	1	2864			
2	8195	1	2870			
2	8196	1	2870			
2	8197	1	2873			
2	8198	1	2873			
2	8199	1	2873			
2	8200	1	2878			
2	8201	1	2878			
2	8202	1	2881			
2	8203	1	2881			
2	8204	1	2884			
2	8205	1	2884			
2	8206	1	2887			
2	8207	1	2887			
2	8208	1	2890			
2	8209	1	2890			
2	8210	1	2893			
2	8211	1	2893			
2	8212	1	2896			
2	8213	1	2896			
2	8214	1	2899			
2	8215	1	2899			
2	8216	1	2902			
2	8217	1	2902			
2	8218	1	2905			
2	8219	1	2905			
2	8220	1	2908			
2	8221	1	2908			
2	8222	1	2908			
2	8223	1	2914			
2	8224	1	2914			
2	8225	1	2917			
2	8226	1	2917			
2	8227	1	2917			
2	8228	1	2923			
2	8229	1	2923			
2	8230	1	2926			
2	8231	1	2926			
2	8232	1	2926			
2	8233	1	2930			
2	8234	1	2930			
2	8235	1	2930			
2	8236	1	2934			
2	8237	1	2934			
2	8238	1	2934			
2	8239	1	2938			
2	8240	1	2938			
2	8241	1	2938			
2	8242	1	2942			
2	8243	1	2942			
2	8244	1	2942			
2	8245	1	2946			
2	8246	1	2946			
2	8247	1	2946			
2	8248	1	2950			
2	8249	1	2950			
2	8250	1	2950			
2	8251	1	2954			
2	8252	1	2954			
2	8253	1	2954			
2	8254	1	2958			
2	8255	1	2958			
2	8256	1	2958			
2	8257	1	2962			
2	8258	1	2962			
2	8259	1	2962			
2	8260	1	2968			
2	8261	1	2968			
2	8262	1	2971			
2	8263	1	2971			
2	8264	1	2971			
2	8265	1	2977			
2	8266	1	2977			
2	8267	1	2980			
2	8268	1	2980			
2	8269	1	2983			
2	8270	1	2983			
2	8271	1	2983			
2	8272	1	3007			
2	8273	1	3007			
2	8274	1	3010			
2	8275	1	3010			
2	8276	1	3010			
2	8277	1	3016			
2	8278	1	3016			
2	8279	1	3019			
2	8280	1	3019			
2	8281	1	3022			
2	8282	1	3022			
2	8283	1	3022			
2	8284	1	3028			
2	8285	1	3028			
2	8286	1	3031			
2	8287	1	3031			
2	8288	1	3034			
2	8289	1	3034			
2	8290	1	3037			
2	8291	1	3037			
2	8292	1	3040			
2	8293	1	3040			
2	8294	1	3043			
2	8295	1	3043			
2	8296	1	3046			
2	8297	1	3046			
2	8298	1	3049			
2	8299	1	3049			
2	8300	1	3052			
2	8301	1	3052			
2	8302	1	3055			
2	8303	1	3055			
2	8304	1	3058			
2	8305	1	3058			
2	8306	1	3058			
2	8307	1	3064			
2	8308	1	3064			
2	8309	1	3067			
2	8310	1	3067			
2	8311	1	3070			
2	8312	1	3070			
2	8313	1	3070			
2	8314	1	3076			
2	8315	1	3076			
2	8316	1	3079			
2	8317	1	3079			
2	8318	1	3079			
2	8319	1	3083			
2	8320	1	3083			
2	8321	1	3083			
2	8322	1	3087			
2	8323	1	3087			
2	8324	1	3087			
2	8325	1	3091			
2	8326	1	3091			
2	8327	1	3091			
2	8328	1	3095			
2	8329	1	3095			
2	8330	1	3095			
2	8331	1	3099			
2	8332	1	3099			
2	8333	1	3099			
2	8334	1	3103			
2	8335	1	3103			
2	8336	1	3103			
2	8337	1	3107			
2	8338	1	3107			
2	8339	1	3107			
2	8340	1	3111			
2	8341	1	3111			
2	8342	1	3111			
2	8343	1	3115			
2	8344	1	3115			
2	8345	1	3115			
2	8346	1	3121			
2	8347	1	3121			
2	8348	1	3124			
2	8349	1	3124			
2	8350	1	3127			
2	8351	1	3127			
2	8352	1	3127			
2	8353	1	3133			
2	8354	1	3133			
2	8355	1	3136			
2	8356	1	3136			
2	8357	1	3136			
2	8358	1	3142			
2	8359	1	3142			
2	8360	1	3147			
2	8361	1	3147			
2	8362	1	3152			
2	8363	1	3152			
2	8364	1	3157			
2	8365	1	3157			
2	8366	1	3162			
2	8367	1	3162			
2	8368	1	3167			
2	8369	1	3167			
2	8370	1	3172			
2	8371	1	3172			
2	8372	1	3177			
2	8373	1	3177			
2	8374	1	3182			
2	8375	1	3182			
2	8376	1	3187			
2	8377	1	3187			
2	8378	1	3190			
2	8379	1	3190			
2	8380	1	3193			
2	8381	1	3193			
2	8382	1	3193			
2	8383	1	3199			
2	8384	1	3199			
2	8385	1	3202			
2	8386	1	3202			
2	8387	1	3202			
2	8388	1	3208			
2	8389	1	3208			
2	8390	1	3212			
2	8391	1	3212			
2	8392	1	3215			
2	8393	1	3215			
2	8394	1	3218			
2	8395	1	3218			
2	8396	1	3221			
2	8397	1	3221			
2	8398	1	3224			
2	8399	1	3224			
2	8400	1	3227			
2	8401	1	3227			
2	8402	1	3230			
2	8403	1	3230			
2	8404	1	3233			
2	8405	1	3233			
2	8406	1	3236			
2	8407	1	3236			
2	8408	1	3239			
2	8409	1	3239			
2	8410	1	3239			
2	8411	1	3245			
2	8412	1	3245			
2	8413	1	3248			
2	8414	1	3248			
2	8415	1	3248			
2	8416	1	3254			
2	8417	1	3254			
2	8418	1	3257			
2	8419	1	3257			
2	8420	1	3260			
2	8421	1	3260			
2	8422	1	3260			
2	8423	1	3264			
2	8424	1	3264			
2	8425	1	3264			
2	8426	1	3268			
2	8427	1	3268			
2	8428	1	3268			
2	8429	1	3272			
2	8430	1	3272			
2	8431	1	3272			
2	8432	1	3276			
2	8433	1	3276			
2	8434	1	3276			
2	8435	1	3280			
2	8436	1	3280			
2	8437	1	3280			
2	8438	1	3284			
2	8439	1	3284			
2	8440	1	3284			
2	8441	1	3288			
2	8442	1	3288			
2	8443	1	3288			
2	8444	1	3292			
2	8445	1	3292			
2	8446	1	3292			
2	8447	1	3296			
2	8448	1	3296			
2	8449	1	3296			
2	8450	1	3302			
2	8451	1	3302			
2	8452	1	3305			
2	8453	1	3305			
2	8454	1	3305			
2	8455	1	3311			
2	8456	1	3311			
2	8457	1	3314			
2	8458	1	3314			
2	8459	1	3317			
2	8460	1	3317			
2	8461	1	3317			
2	8462	1	3341			
2	8463	1	3341			
2	8464	1	3344			
2	8465	1	3344			
2	8466	1	3344			
2	8467	1	3350			
2	8468	1	3350			
2	8469	1	3353			
2	8470	1	3353			
2	8471	1	3356			
2	8472	1	3356			
2	8473	1	3356			
2	8474	1	3362			
2	8475	1	3362			
2	8476	1	3365			
2	8477	1	3365			
2	8478	1	3368			
2	8479	1	3368			
2	8480	1	3371			
2	8481	1	3371			
2	8482	1	3374			
2	8483	1	3374			
2	8484	1	3377			
2	8485	1	3377			
2	8486	1	3380			
2	8487	1	3380			
2	8488	1	3383			
2	8489	1	3383			
2	8490	1	3386			
2	8491	1	3386			
2	8492	1	3389			
2	8493	1	3389			
2	8494	1	3392			
2	8495	1	3392			
2	8496	1	3392			
2	8497	1	3398			
2	8498	1	3398			
2	8499	1	3401			
2	8500	1	3401			
2	8501	1	3404			
2	8502	1	3404			
2	8503	1	3404			
2	8504	1	3410			
2	8505	1	3410			
2	8506	1	3413			
2	8507	1	3413			
2	8508	1	3413			
2	8509	1	3417			
2	8510	1	3417			
2	8511	1	3417			
2	8512	1	3421			
2	8513	1	3421			
2	8514	1	3421			
2	8515	1	3425			
2	8516	1	3425			
2	8517	1	3425			
2	8518	1	3429			
2	8519	1	3429			
2	8520	1	3429			
2	8521	1	3433			
2	8522	1	3433			
2	8523	1	3433			
2	8524	1	3437			
2	8525	1	3437			
2	8526	1	3437			
2	8527	1	3441			
2	8528	1	3441			
2	8529	1	3441			
2	8530	1	3445			
2	8531	1	3445			
2	8532	1	3445			
2	8533	1	3449			
2	8534	1	3449			
2	8535	1	3449			
2	8536	1	3455			
2	8537	1	3455			
2	8538	1	3458			
2	8539	1	3458			
2	8540	1	3461			
2	8541	1	3461			
2	8542	1	3461			
2	8543	1	3467			
2	8544	1	3467			
2	8545	1	3470			
2	8546	1	3470			
2	8547	1	3470			
2	8548	1	3476			
2	8549	1	3476			
2	8550	1	3481			
2	8551	1	3481			
2	8552	1	3486			
2	8553	1	3486			
2	8554	1	3491			
2	8555	1	3491			
2	8556	1	3496			
2	8557	1	3496			
2	8558	1	3501			
2	8559	1	3501			
2	8560	1	3506			
2	8561	1	3506			
2	8562	1	3511			
2	8563	1	3511			
2	8564	1	3516			
2	8565	1	3516			
2	8566	1	3521			
2	8567	1	3521			
2	8568	1	3524			
2	8569	1	3524			
2	8570	1	3527			
2	8571	1	3527			
2	8572	1	3527			
2	8573	1	3533			
2	8574	1	3533			
2	8575	1	3536			
2	8576	1	3536			
2	8577	1	3536			
2	8578	1	3542			
2	8579	1	3542			
2	8580	1	3545			
2	8581	1	3545			
2	8582	1	3548			
2	8583	1	3548			
2	8584	1	3548			
2	8585	1	3553			
2	8586	1	3553			
2	8587	1	3556			
2	8588	1	3556			
2	8589	1	3559			
2	8590	1	3559			
2	8591	1	3562			
2	8592	1	3562			
2	8593	1	3565			
2	8594	1	3565			
2	8595	1	3568			
2	8596	1	3568			
2	8597	1	3571			
2	8598	1	3571			
2	8599	1	3574			
2	8600	1	3574			
2	8601	1	3577			
2	8602	1	3577			
2	8603	1	3577			
2	8604	1	3583			
2	8605	1	3583			
2	8606	1	3586			
2	8607	1	3586			
2	8608	1	3586			
2	8609	1	3592			
2	8610	1	3592			
2	8611	1	3595			
2	8612	1	3595			
2	8613	1	3598			
2	8614	1	3598			
2	8615	1	3598			
2	8616	1	3604			
2	8617	1	3604			
2	8618	1	3604			
2	8619	1	3608			
2	8620	1	3608			
2	8621	1	3608			
2	8622	1	3612			
2	8623	1	3612			
2	8624	1	3612			
2	8625	1	3616			
2	8626	1	3616			
2	8627	1	3616			
2	8628	1	3620			
2	8629	1	3620			
2	8630	1	3620			
2	8631	1	3624			
2	8632	1	3624			
2	8633	1	3624			
2	8634	1	3628			
2	8635	1	3628			
2	8636	1	3628			
2	8637	1	3632			
2	8638	1	3632			
2	8639	1	3632			
2	8640	1	3638			
2	8641	1	3638			
2	8642	1	3641			
2	8643	1	3641			
2	8644	1	3641			
2	8645	1	3647			
2	8646	1	3647			
2	8647	1	3650			
2	8648	1	3650			
2	8649	1	3653			
2	8650	1	3653			
2	8651	1	3653			
2	8652	1	3659			
2	8653	1	3659			
2	8654	1	3678			
2	8655	1	3678			
2	8656	1	3681			
2	8657	1	3681			
2	8658	1	3681			
2	8659	1	3687			
2	8660	1	3687			
2	8661	1	3690			
2	8662	1	3690			
2	8663	1	3693			
2	8664	1	3693			
2	8665	1	3693			
2	8666	1	3699			
2	8667	1	3699			
2	8668	1	3702			
2	8669	1	3702			
2	8670	1	3702			
2	8671	1	3706			
2	8672	1	3706			
2	8673	1	3709			
2	8674	1	3709			
2	8675	1	3712			
2	8676	1	3712			
2	8677	1	3715			
2	8678	1	3715			
2	8679	1	3718			
2	8680	1	3718			
2	8681	1	3721			
2	8682	1	3721			
2	8683	1	3724			
2	8684	1	3724			
2	8685	1	3727			
2	8686	1	3727			
2	8687	1	3730			
2	8688	1	3730			
2	8689	1	3730			
2	8690	1	3736			
2	8691	1	3736			
2	8692	1	3739			
2	8693	1	3739			
2	8694	1	3742			
2	8695	1	3742			
2	8696	1	3742			
2	8697	1	3748			
2	8698	1	3748			
2	8699	1	3751			
2	8700	1	3751			
2	8701	1	3751			
2	8702	1	3757			
2	8703	1	3757			
2	8704	1	3760			
2	8705	1	3760			
2	8706	1	3760			
2	8707	1	3764			
2	8708	1	3764			
2	8709	1	3764			
2	8710	1	3768			
2	8711	1	3768			
2	8712	1	3768			
2	8713	1	3772			
2	8714	1	3772			
2	8715	1	3772			
2	8716	1	3776			
2	8717	1	3776			
2	8718	1	3776			
2	8719	1	3780			
2	8720	1	3780			
2	8721	1	3780			
2	8722	1	3784			
2	8723	1	3784			
2	8724	1	3784			
2	8725	1	3788			
2	8726	1	3788			
2	8727	1	3788			
2	8728	1	3794			
2	8729	1	3794			
2	8730	1	3797			
2	8731	1	3797			
2	8732	1	3800			
2	8733	1	3800			
2	8734	1	3800			
2	8735	1	3806			
2	8736	1	3806			
2	8737	1	3809			
2	8738	1	3809			
2	8739	1	3809			
2	8740	1	3815			
2	8741	1	3815			
2	8742	1	3818			
2	8743	1	3818			
2	8744	1	3821			
2	8745	1	3821			
2	8746	1	3821			
2	8747	1	3827			
2	8748	1	3827			
2	8749	1	3832			
2	8750	1	3832			
2	8751	1	3837			
2	8752	1	3837			
2	8753	1	3842			
2	8754	1	3842			
2	8755	1	3847			
2	8756	1	3847			
2	8757	1	3852			
2	8758	1	3852			
2	8759	1	3857			
2	8760	1	3857			
2	8761	1	3862			
2	8762	1	3862			
2	8763	1	3865			
2	8764	1	3865			
2	8765	1	3868			
2	8766	1	3868			
2	8767	1	3868			
2	8768	1	3874			
2	8769	1	3874			
2	8770	1	3877			
2	8771	1	3877			
2	8772	1	3877			
2	8773	1	3883			
2	8774	1	3883			
2	8775	1	3886			
2	8776	1	3886			
2	8777	1	3889			
2	8778	1	3889			
2	8779	1	3889			
2	8780	1	3896			
2	8781	1	3896			
2	8782	1	3899			
2	8783	1	3899			
2	8784	1	3902			
2	8785	1	3902			
2	8786	1	3905			
2	8787	1	3905			
2	8788	1	3908			
2	8789	1	3908			
2	8790	1	3911			
2	8791	1	3911			
2	8792	1	3914			
2	8793	1	3914			
2	8794	1	3917			
2	8795	1	3917			
2	8796	1	3917			
2	8797	1	3923			
2	8798	1	3923			
2	8799	1	3926			
2	8800	1	3926			
2	8801	1	3926			
2	8802	1	3932			
2	8803	1	3932			
2	8804	1	3935			
2	8805	1	3935			
2	8806	1	3938			
2	8807	1	3938			
2	8808	1	3938			
2	8809	1	3944			
2	8810	1	3944			
2	8811	1	3947			
2	8812	1	3947			
2	8813	1	3947			
2	8814	1	3951			
2	8815	1	3951			
2	8816	1	3951			
2	8817	1	3955			
2	8818	1	3955			
2	8819	1	3955			
2	8820	1	3959			
2	8821	1	3959			
2	8822	1	3959			
2	8823	1	3963			
2	8824	1	3963			
2	8825	1	3963			
2	8826	1	3967			
2	8827	1	3967			
2	8828	1	3967			
2	8829	1	3971			
2	8830	1	3971			
2	8831	1	3971			
2	8832	1	3977			
2	8833	1	3977			
2	8834	1	3980			
2	8835	1	3980			
2	8836	1	3980			
2	8837	1	3986			
2	8838	1	3986			
2	8839	1	3989			
2	8840	1	3989			
2	8841	1	3992			
2	8842	1	3992			
2	8843	1	3992			
2	8844	1	3998			
2	8845	1	3998			
2	8846	1	4001			
2	8847	1	4001			
2	8848	1	4001			
2	8849	1	4019			
2	8850	1	4019			
2	8851	1	4022			
2	8852	1	4022			
2	8853	1	4022			
2	8854	1	4028			
2	8855	1	4028			
2	8856	1	4031			
2	8857	1	4031			
2	8858	1	4034			
2	8859	1	4034			
2	8860	1	4034			
2	8861	1	4040			
2	8862	1	4040			
2	8863	1	4043			
2	8864	1	4043			
2	8865	1	4043			
2	8866	1	4049			
2	8867	1	4049			
2	8868	1	4052			
2	8869	1	4052			
2	8870	1	4055			
2	8871	1	4055			
2	8872	1	4058			
2	8873	1	4058			
2	8874	1	4061			
2	8875	1	4061			
2	8876	1	4064			
2	8877	1	4064			
2	8878	1	4067			
2	8879	1	4067			
2	8880	1	4070			
2	8881	1	4070			
2	8882	1	4073			
2	8883	1	4073			
2	8884	1	4073			
2	8885	1	4079			
2	8886	1	4079			
2	8887	1	4082			
2	8888	1	4082			
2	8889	1	4085			
2	8890	1	4085			
2	8891	1	4085			
2	8892	1	4091			
2	8893	1	4091			
2	8894	1	4094			
2	8895	1	4094			
2	8896	1	4094			
2	8897	1	4100			
2	8898	1	4100			
2	8899	1	4103			
2	8900	1	4103			
2	8901	1	4106			
2	8902	1	4106			
2	8903	1	4106			
2	8904	1	4110			
2	8905	1	4110			
2	8906	1	4110			
2	8907	1	4114			
2	8908	1	4114			
2	8909	1	4114			
2	8910	1	4118			
2	8911	1	4118			
2	8912	1	4118			
2	8913	1	4122			
2	8914	1	4122			
2	8915	1	4122			
2	8916	1	4126			
2	8917	1	4126			
2	8918	1	4126			
2	8919	1	4130			
2	8920	1	4130			
2	8921	1	4130			
2	8922	1	4134			
2	8923	1	4134			
2	8924	1	4134			
2	8925	1	4140			
2	8926	1	4140			
2	8927	1	4143			
2	8928	1	4143			
2	8929	1	4146			
2	8930	1	4146			
2	8931	1	4146			
2	8932	1	4152			
2	8933	1	4152			
2	8934	1	4155			
2	8935	1	4155			
2	8936	1	4155			
2	8937	1	4161			
2	8938	1	4161			
2	8939	1	4164			
2	8940	1	4164			
2	8941	1	4167			
2	8942	1	4167			
2	8943	1	4167			
2	8944	1	4175			
2	8945	1	4175			
2	8946	1	4180			
2	8947	1	4180			
2	8948	1	4185			
2	8949	1	4185			
2	8950	1	4190			
2	8951	1	4190			
2	8952	1	4195			
2	8953	1	4195			
2	8954	1	4200			
2	8955	1	4200			
2	8956	1	4205			
2	8957	1	4205			
2	8958	1	4208			
2	8959	1	4208			
2	8960	1	4211			
2	8961	1	4211			
2	8962	1	4211			
2	8963	1	4217			
2	8964	1	4217			
2	8965	1	4220			
2	8966	1	4220			
2	8967	1	4220			
2	8968	1	4226			
2	8969	1	4226			
2	8970	1	4229			
2	8971	1	4229			
2	8972	1	4232			
2	8973	1	4232			
2	8974	1	4232			
2	8975	1	4238			
2	8976	1	4238			
2	8977	1	4242			
2	8978	1	4242			
2	8979	1	4245			
2	8980	1	4245			
2	8981	1	4248			
2	8982	1	4248			
2	8983	1	4251			
2	8984	1	4251			
2	8985	1	4254			
2	8986	1	4254			
2	8987	1	4257			
2	8988	1	4257			
2	8989	1	4260			
2	8990	1	4260			
2	8991	1	4260			
2	8992	1	4266			
2	8993	1	4266			
2	8994	1	4269			
2	8995	1	4269			
2	8996	1	4269			
2	8997	1	4275			
2	8998	1	4275			
2	8999	1	4278			
2	9000	1	4278			
2	9001	1	4281			
2	9002	1	4281			
2	9003	1	4281			
2	9004	1	4287			
2	9005	1	4287			
2	9006	1	4290			
2	9007	1	4290			
2	9008	1	4290			
2	9009	1	4294			
2	9010	1	4294			
2	9011	1	4294			
2	9012	1	4298			
2	9013	1	4298			
2	9014	1	4298			
2	9015	1	4302			
2	9016	1	4302			
2	9017	1	4302			
2	9018	1	4306			
2	9019	1	4306			
2	9020	1	4306			
2	9021	1	4310			
2	9022	1	4310			
2	9023	1	4310			
2	9024	1	4314			
2	9025	1	4314			
2	9026	1	4314			
2	9027	1	4320			
2	9028	1	4320			
2	9029	1	4323			
2	9030	1	4323			
2	9031	1	4323			
2	9032	1	4329			
2	9033	1	4329			
2	9034	1	4332			
2	9035	1	4332			
2	9036	1	4335			
2	9037	1	4335			
2	9038	1	4335			
2	9039	1	4341			
2	9040	1	4341			
2	9041	1	4344			
2	9042	1	4344			
2	9043	1	4344			
2	9044	1	4350			
2	9045	1	4350			
2	9046	1	4365			
2	9047	1	4365			
2	9048	1	4368			
2	9049	1	4368			
2	9050	1	4368			
2	9051	1	4374			
2	9052	1	4374			
2	9053	1	4377			
2	9054	1	4377			
2	9055	1	4380			
2	9056	1	4380			
2	9057	1	4380			
2	9058	1	4386			
2	9059	1	4386			
2	9060	1	4389			
2	9061	1	4389			
2	9062	1	4389			
2	9063	1	4395			
2	9064	1	4395			
2	9065	1	4398			
2	9066	1	4398			
2	9067	1	4401			
2	9068	1	4401			
2	9069	1	4401			
2	9070	1	4405			
2	9071	1	4405			
2	9072	1	4408			
2	9073	1	4408			
2	9074	1	4411			
2	9075	1	4411			
2	9076	1	4414			
2	9077	1	4414			
2	9078	1	4417			
2	9079	1	4417			
2	9080	1	4420			
2	9081	1	4420			
2	9082	1	4423			
2	9083	1	4423			
2	9084	1	4423			
2	9085	1	4429			
2	9086	1	4429			
2	9087	1	4432			
2	9088	1	4432			
2	9089	1	4435			
2	9090	1	4435			
2	9091	1	4435			
2	9092	1	4441			
2	9093	1	4441			
2	9094	1	4444			
2	9095	1	4444			
2	9096	1	4444			
2	9097	1	4450			
2	9098	1	4450			
2	9099	1	4453			
2	9100	1	4453			
2	9101	1	4456			
2	9102	1	4456			
2	9103	1	4456			
2	9104	1	4462			
2	9105	1	4462			
2	9106	1	4462			
2	9107	1	4466			
2	9108	1	4466			
2	9109	1	4466			
2	9110	1	4470			
2	9111	1	4470			
2	9112	1	4470			
2	9113	1	4474			
2	9114	1	4474			
2	9115	1	4474			
2	9116	1	4478			
2	9117	1	4478			
2	9118	1	4478			
2	9119	1	4482			
2	9120	1	4482			
2	9121	1	4482			
2	9122	1	4488			
2	9123	1	4488			
2	9124	1	4491			
2	9125	1	4491			
2	9126	1	4494			
2	9127	1	4494			
2	9128	1	4494			
2	9129	1	4500			
2	9130	1	4500			
2	9131	1	4503			
2	9132	1	4503			
2	9133	1	4503			
2	9134	1	4509			
2	9135	1	4509			
2	9136	1	4512			
2	9137	1	4512			
2	9138	1	4515			
2	9139	1	4515			
2	9140	1	4515			
2	9141	1	4521			
2	9142	1	4521			
2	9143	1	4526			
2	9144	1	4526			
2	9145	1	4531			
2	9146	1	4531			
2	9147	1	4536			
2	9148	1	4536			
2	9149	1	4541			
2	9150	1	4541			
2	9151	1	4546			
2	9152	1	4546			
2	9153	1	4551			
2	9154	1	4551			
2	9155	1	4554			
2	9156	1	4554			
2	9157	1	4557			
2	9158	1	4557			
2	9159	1	4557			
2	9160	1	4563			
2	9161	1	4563			
2	9162	1	4566			
2	9163	1	4566			
2	9164	1	4566			
2	9165	1	4572			
2	9166	1	4572			
2	9167	1	4575			
2	9168	1	4575			
2	9169	1	4578			
2	9170	1	4578			
2	9171	1	4578			
2	9172	1	4584			
2	9173	1	4584			
2	9174	1	4587			
2	9175	1	4587			
2	9176	1	4587			
2	9177	1	4592			
2	9178	1	4592			
2	9179	1	4595			
2	9180	1	4595			
2	9181	1	4598			
2	9182	1	4598			
2	9183	1	4601			
2	9184	1	4601			
2	9185	1	4604			
2	9186	1	4604			
2	9187	1	4607			
2	9188	1	4607			
2	9189	1	4607			
2	9190	1	4613			
2	9191	1	4613			
2	9192	1	4616			
2	9193	1	4616			
2	9194	1	4616			
2	9195	1	4622			
2	9196	1	4622			
2	9197	1	4625			
2	9198	1	4625			
2	9199	1	4628			
2	9200	1	4628			
2	9201	1	4628			
2	9202	1	4634			
2	9203	1	4634			
2	9204	1	4637			
2	9205	1	4637			
2	9206	1	4637			
2	9207	1	4643			
2	9208	1	4643			
2	9209	1	4646			
2	9210	1	4646			
2	9211	1	4646			
2	9212	1	4650			
2	9213	1	4650			
2	9214	1	4650			
2	9215	1	4654			
2	9216	1	4654			
2	9217	1	4654			
2	9218	1	4658			
2	9219	1	4658			
2	9220	1	4658			
2	9221	1	4662			
2	9222	1	4662			
2	9223	1	4662			
2	9224	1	4668			
2	9225	1	4668			
2	9226	1	4671			
2	9227	1	4671			
2	9228	1	4671			
2	9229	1	4677			
2	9230	1	4677			
2	9231	1	4680			
2	9232	1	4680			
2	9233	1	4683			
2	9234	1	4683			
2	9235	1	4683			
2	9236	1	4689			
2	9237	1	4689			
2	9238	1	4692			
2	9239	1	4692			
2	9240	1	4692			
2	9241	1	4698			
2	9242	1	4698			
2	9243	1	4701			
2	9244	1	4701			
2	9245	1	4704			
2	9246	1	4704			
2	9247	1	4704			
2	9248	1	4718			
2	9249	1	4718			
2	9250	1	4721			
2	9251	1	4721			
2	9252	1	4721			
2	9253	1	4727			
2	9254	1	4727			
2	9255	1	4730			
2	9256	1	4730			
2	9257	1	4733			
2	9258	1	4733			
2	9259	1	4733			
2	9260	1	4739			
2	9261	1	4739			
2	9262	1	4742			
2	9263	1	4742			
2	9264	1	4742			
2	9265	1	4748			
2	9266	1	4748			
2	9267	1	4751			
2	9268	1	4751			
2	9269	1	4754			
2	9270	1	4754			
2	9271	1	4754			
2	9272	1	4760			
2	9273	1	4760			
2	9274	1	4763			
2	9275	1	4763			
2	9276	1	4766			
2	9277	1	4766			
2	9278	1	4769			
2	9279	1	4769			
2	9280	1	4772			
2	9281	1	4772			
2	9282	1	4775			
2	9283	1	4775			
2	9284	1	4775			
2	9285	1	4781			
2	9286	1	4781			
2	9287	1	4784			
2	9288	1	4784			
2	9289	1	4787			
2	9290	1	4787			
2	9291	1	4787			
2	9292	1	4793			
2	9293	1	4793			
2	9294	1	4796			
2	9295	1	4796			
2	9296	1	4796			
2	9297	1	4802			
2	9298	1	4802			
2	9299	1	4805			
2	9300	1	4805			
2	9301	1	4808			
2	9302	1	4808			
2	9303	1	4808			
2	9304	1	4814			
2	9305	1	4814			
2	9306	1	4817			
2	9307	1	4817			
2	9308	1	4817			
2	9309	1	4821			
2	9310	1	4821			
2	9311	1	4821			
2	9312	1	4825			
2	9313	1	4825			
2	9314	1	4825			
2	9315	1	4829			
2	9316	1	4829			
2	9317	1	4829			
2	9318	1	4833			
2	9319	1	4833			
2	9320	1	4833			
2	9321	1	4839			
2	9322	1	4839			
2	9323	1	4842			
2	9324	1	4842			
2	9325	1	4845			
2	9326	1	4845			
2	9327	1	4845			
2	9328	1	4851			
2	9329	1	4851			
2	9330	1	4854			
2	9331	1	4854			
2	9332	1	4854			
2	9333	1	4860			
2	9334	1	4860			
2	9335	1	4863			
2	9336	1	4863			
2	9337	1	4866			
2	9338	1	4866			
2	9339	1	4866			
2	9340	1	4872			
2	9341	1	4872			
2	9342	1	4875			
2	9343	1	4875			
2	9344	1	4875			
2	9345	1	4881			
2	9346	1	4881			
2	9347	1	4886			
2	9348	1	4886			
2	9349	1	4891			
2	9350	1	4891			
2	9351	1	4896			
2	9352	1	4896			
2	9353	1	4901			
2	9354	1	4901			
2	9355	1	4904			
2	9356	1	4904			
2	9357	1	4907			
2	9358	1	4907			
2	9359	1	4907			
2	9360	1	4913			
2	9361	1	4913			
2	9362	1	4916			
2	9363	1	4916			
2	9364	1	4916			
2	9365	1	4922			
2	9366	1	4922			
2	9367	1	4925			
2	9368	1	4925			
2	9369	1	4928			
2	9370	1	4928			
2	9371	1	4928			
2	9372	1	4934			
2	9373	1	4934			
2	9374	1	4937			
2	9375	1	4937			
2	9376	1	4937			
2	9377	1	4943			
2	9378	1	4943			
2	9379	1	4947			
2	9380	1	4947			
2	9381	1	4950			
2	9382	1	4950			
2	9383	1	4953			
2	9384	1	4953			
2	9385	1	4956			
2	9386	1	4956			
2	9387	1	4959			
2	9388	1	4959			
2	9389	1	4959			
2	9390	1	4965			
2	9391	1	4965			
2	9392	1	4968			
2	9393	1	4968			
2	9394	1	4968			
2	9395	1	4974			
2	9396	1	4974			
2	9397	1	4977			
2	9398	1	4977			
2	9399	1	4980			
2	9400	1	4980			
2	9401	1	4980			
2	9402	1	4986			
2	9403	1	4986			
2	9404	1	4989			
2	9405	1	4989			
2	9406	1	4989			
2	9407	1	4995			
2	9408	1	4995			
2	9409	1	4998			
2	9410	1	4998			
2	9411	1	5001			
2	9412	1	5001			
2	9413	1	5001			
2	9414	1	5005			
2	9415	1	5005			
2	9416	1	5005			
2	9417	1	5009			
2	9418	1	5009			
2	9419	1	5009			
2	9420	1	5013			
2	9421	1	5013			
2	9422	1	5013			
2	9423	1	5017			
2	9424	1	5017			
2	9425	1	5017			
2	9426	1	5023			
2	9427	1	5023			
2	9428	1	5026			
2	9429	1	5026			
2	9430	1	5026			
2	9431	1	5032			
2	9432	1	5032			
2	9433	1	5035			
2	9434	1	5035			
2	9435	1	5038			
2	9436	1	5038			
2	9437	1	5038			
2	9438	1	5044			
2	9439	1	5044			
2	9440	1	5047			
2	9441	1	5047			
2	9442	1	5047			
2	9443	1	5053			
2	9444	1	5053			
2	9445	1	5056			
2	9446	1	5056			
2	9447	1	5059			
2	9448	1	5059			
2	9449	1	5059			
2	9450	1	5073			
2	9451	1	5073			
2	9452	1	5076			
2	9453	1	5076			
2	9454	1	5076			
2	9455	1	5082			
2	9456	1	5082			
2	9457	1	5085			
2	9458	1	5085			
2	9459	1	5088			
2	9460	1	5088			
2	9461	1	5088			
2	9462	1	5094			
2	9463	1	5094			
2	9464	1	5097			
2	9465	1	5097			
2	9466	1	5097			
2	9467	1	5103			
2	9468	1	5103			
2	9469	1	5106			
2	9470	1	5106			
2	9471	1	5109			
2	9472	1	5109			
2	9473	1	5109			
2	9474	1	5115			
2	9475	1	5115			
2	9476	1	5118			
2	9477	1	5118			
2	9478	1	5121			
2	9479	1	5121			
2	9480	1	5124			
2	9481	1	5124			
2	9482	1	5127			
2	9483	1	5127			
2	9484	1	5130			
2	9485	1	5130			
2	9486	1	5130			
2	9487	1	5136			
2	9488	1	5136			
2	9489	1	5139			
2	9490	1	5139			
2	9491	1	5142			
2	9492	1	5142			
2	9493	1	5142			
2	9494	1	5148			
2	9495	1	5148			
2	9496	1	5151			
2	9497	1	5151			
2	9498	1	5151			
2	9499	1	5157			
2	9500	1	5157			
2	9501	1	5160			
2	9502	1	5160			
2	9503	1	5163			
2	9504	1	5163			
2	9505	1	5163			
2	9506	1	5169			
2	9507	1	5169			
2	9508	1	5172			
2	9509	1	5172			
2	9510	1	5172			
2	9511	1	5176			
2	9512	1	5176			
2	9513	1	5176			
2	9514	1	5180			
2	9515	1	5180			
2	9516	1	5180			
2	9517	1	5184			
2	9518	1	5184			
2	9519	1	5184			
2	9520	1	5188			
2	9521	1	5188			
2	9522	1	5188			
2	9523	1	5194			
2	9524	1	5194			
2	9525	1	5197			
2	9526	1	5197			
2	9527	1	5200			
2	9528	1	5200			
2	9529	1	5200			
2	9530	1	5206			
2	9531	1	5206			
2	9532	1	5209			
2	9533	1	5209			
2	9534	1	5209			
2	9535	1	5215			
2	9536	1	5215			
2	9537	1	5218			
2	9538	1	5218			
2	9539	1	5221			
2	9540	1	5221			
2	9541	1	5221			
2	9542	1	5227			
2	9543	1	5227			
2	9544	1	5230			
2	9545	1	5230			
2	9546	1	5230			
2	9547	1	5236			
2	9548	1	5236			
2	9549	1	5241			
2	9550	1	5241			
2	9551	1	5246			
2	9552	1	5246			
2	9553	1	5251			
2	9554	1	5251			
2	9555	1	5256			
2	9556	1	5256			
2	9557	1	5259			
2	9558	1	5259			
2	9559	1	5262			
2	9560	1	5262			
2	9561	1	5262			
2	9562	1	5268			
2	9563	1	5268			
2	9564	1	5271			
2	9565	1	5271			
2	9566	1	5271			
2	9567	1	5277			
2	9568	1	5277			
2	9569	1	5280			
2	9570	1	5280			
2	9571	1	5283			
2	9572	1	5283			
2	9573	1	5283			
2	9574	1	5289			
2	9575	1	5289			
2	9576	1	5292			
2	9577	1	5292			
2	9578	1	5292			
2	9579	1	5298			
2	9580	1	5298			
2	9581	1	5301			
2	9582	1	5301			
2	9583	1	5304			
2	9584	1	5304			
2	9585	1	5304			
2	9586	1	5309			
2	9587	1	5309			
2	9588	1	5312			
2	9589	1	5312			
2	9590	1	5315			
2	9591	1	5315			
2	9592	1	5318			
2	9593	1	5318			
2	9594	1	5318			
2	9595	1	5324			
2	9596	1	5324			
2	9597	1	5327			
2	9598	1	5327			
2	9599	1	5327			
2	9600	1	5333			
2	9601	1	5333			
2	9602	1	5336			
2	9603	1	5336			
2	9604	1	5339			
2	9605	1	5339			
2	9606	1	5339			
2	9607	1	5345			
2	9608	1	5345			
2	9609	1	5348			
2	9610	1	5348			
2	9611	1	5348			
2	9612	1	5354			
2	9613	1	5354			
2	9614	1	5357			
2	9615	1	5357			
2	9616	1	5360			
2	9617	1	5360			
2	9618	1	5360			
2	9619	1	5366			
2	9620	1	5366			
2	9621	1	5366			
2	9622	1	5370			
2	9623	1	5370			
2	9624	1	5370			
2	9625	1	5374			
2	9626	1	5374			
2	9627	1	5374			
2	9628	1	5380			
2	9629	1	5380			
2	9630	1	5383			
2	9631	1	5383			
2	9632	1	5383			
2	9633	1	5389			
2	9634	1	5389			
2	9635	1	5392			
2	9636	1	5392			
2	9637	1	5395			
2	9638	1	5395			
2	9639	1	5395			
2	9640	1	5401			
2	9641	1	5401			
2	9642	1	5404			
2	9643	1	5404			
2	9644	1	5404			
2	9645	1	5410			
2	9646	1	5410			
2	9647	1	5413			
2	9648	1	5413			
2	9649	1	5416			
2	9650	1	5416			
2	9651	1	5416			
2	9652	1	5422			
2	9653	1	5422			
2	9654	1	5431			
2	9655	1	5431			
2	9656	1	5434			
2	9657	1	5434			
2	9658	1	5434			
2	9659	1	5440			
2	9660	1	5440			
2	9661	1	5443			
2	9662	1	5443			
2	9663	1	5446			
2	9664	1	5446			
2	9665	1	5446			
2	9666	1	5452			
2	9667	1	5452			
2	9668	1	5455			
2	9669	1	5455			
2	9670	1	5455			
2	9671	1	5461			
2	9672	1	5461			
2	9673	1	5464			
2	9674	1	5464			
2	9675	1	5467			
2	9676	1	5467			
2	9677	1	5467			
2	9678	1	5473			
2	9679	1	5473			
2	9680	1	5476			
2	9681	1	5476			
2	9682	1	5476			
2	9683	1	5480			
2	9684	1	5480			
2	9685	1	5483			
2	9686	1	5483			
2	9687	1	5486			
2	9688	1	5486			
2	9689	1	5489			
2	9690	1	5489			
2	9691	1	5489			
2	9692	1	5495			
2	9693	1	5495			
2	9694	1	5498			
2	9695	1	5498			
2	9696	1	5501			
2	9697	1	5501			
2	9698	1	5501			
2	9699	1	5507			
2	9700	1	5507			
2	9701	1	5510			
2	9702	1	5510			
2	9703	1	5510			
2	9704	1	5516			
2	9705	1	5516			
2	9706	1	5519			
2	9707	1	5519			
2	9708	1	5522			
2	9709	1	5522			
2	9710	1	5522			
2	9711	1	5528			
2	9712	1	5528			
2	9713	1	5531			
2	9714	1	5531			
2	9715	1	5531			
2	9716	1	5537			
2	9717	1	5537			
2	9718	1	5540			
2	9719	1	5540			
2	9720	1	5540			
2	9721	1	5544			
2	9722	1	5544			
2	9723	1	5544			
2	9724	1	5548			
2	9725	1	5548			
2	9726	1	5548			
2	9727	1	5554			
2	9728	1	5554			
2	9729	1	5557			
2	9730	1	5557			
2	9731	1	5560			
2	9732	1	5560			
2	9733	1	5560			
2	9734	1	5566			
2	9735	1	5566			
2	9736	1	5569			
2	9737	1	5569			
2	9738	1	5569			
2	9739	1	5575			
2	9740	1	5575			
2	9741	1	5578			
2	9742	1	5578			
2	9743	1	5581			
2	9744	1	5581			
2	9745	1	5581			
2	9746	1	5587			
2	9747	1	5587			
2	9748	1	5590			
2	9749	1	5590			
2	9750	1	5590			
2	9751	1	5596			
2	9752	1	5596			
2	9753	1	5599			
2	9754	1	5599			
2	9755	1	5602			
2	9756	1	5602			
2	9757	1	5602			
2	9758	1	5608			
2	9759	1	5608			
2	9760	1	5613			
2	9761	1	5613			
2	9762	1	5618			
2	9763	1	5618			
2	9764	1	5621			
2	9765	1	5621			
2	9766	1	5624			
2	9767	1	5624			
2	9768	1	5624			
2	9769	1	5630			
2	9770	1	5630			
2	9771	1	5633			
2	9772	1	5633			
2	9773	1	5633			
2	9774	1	5639			
2	9775	1	5639			
2	9776	1	5642			
2	9777	1	5642			
2	9778	1	5645			
2	9779	1	5645			
2	9780	1	5645			
2	9781	1	5651			
2	9782	1	5651			
2	9783	1	5654			
2	9784	1	5654			
2	9785	1	5654			
2	9786	1	5660			
2	9787	1	5660			
2	9788	1	5663			
2	9789	1	5663			
2	9790	1	5666			
2	9791	1	5666			
2	9792	1	5666			
2	9793	1	5673			
2	9794	1	5673			
2	9795	1	5676			
2	9796	1	5676			
2	9797	1	5679			
2	9798	1	5679			
2	9799	1	5679			
2	9800	1	5685			
2	9801	1	5685			
2	9802	1	5688			
2	9803	1	5688			
2	9804	1	5688			
2	9805	1	5694			
2	9806	1	5694			
2	9807	1	5697			
2	9808	1	5697			
2	9809	1	5700			
2	9810	1	5700			
2	9811	1	5700			
2	9812	1	5706			
2	9813	1	5706			
2	9814	1	5709			
2	9815	1	5709			
2	9816	1	5709			
2	9817	1	5715			
2	9818	1	5715			
2	9819	1	5718			
2	9820	1	5718			
2	9821	1	5721			
2	9822	1	5721			
2	9823	1	5721			
2	9824	1	5727			
2	9825	1	5727			
2	9826	1	5730			
2	9827	1	5730			
2	9828	1	5730			
2	9829	1	5734			
2	9830	1	5734			
2	9831	1	5734			
2	9832	1	5740			
2	9833	1	5740			
2	9834	1	5743			
2	9835	1	5743			
2	9836	1	5743			
2	9837	1	5749			
2	9838	1	5749			
2	9839	1	5752			
2	9840	1	5752			
2	9841	1	5755			
2	9842	1	5755			
2	9843	1	5755			
2	9844	1	5761			
2	9845	1	5761			
2	9846	1	5764			
2	9847	1	5764			
2	9848	1	5764			
2	9849	1	5770			
2	9850	1	5770			
2	9851	1	5773			
2	9852	1	5773			
2	9853	1	5776			
2	9854	1	5776			
2	9855	1	5776			
2	9856	1	5782			
2	9857	1	5782			
2	9858	1	5789			
2	9859	1	5789			
2	9860	1	5792			
2	9861	1	5792			
2	9862	1	5792			
2	9863	1	5798			
2	9864	1	5798			
2	9865	1	5801			
2	9866	1	5801			
2	9867	1	5804			
2	9868	1	5804			
2	9869	1	5804			
2	9870	1	5810			
2	9871	1	5810			
2	9872	1	5813			
2	9873	1	5813			
2	9874	1	5813			
2	9875	1	5819			
2	9876	1	5819			
2	9877	1	5822			
2	9878	1	5822			
2	9879	1	5825			
2	9880	1	5825			
2	9881	1	5825			
2	9882	1	5831			
2	9883	1	5831			
2	9884	1	5834			
2	9885	1	5834			
2	9886	1	5837			
2	9887	1	5837			
2	9888	1	5840			
2	9889	1	5840			
2	9890	1	5840			
2	9891	1	5846			
2	9892	1	5846			
2	9893	1	5849			
2	9894	1	5849			
2	9895	1	5852			
2	9896	1	5852			
2	9897	1	5852			
2	9898	1	5858			
2	9899	1	5858			
2	9900	1	5861			
2	9901	1	5861			
2	9902	1	5861			
2	9903	1	5867			
2	9904	1	5867			
2	9905	1	5870			
2	9906	1	5870			
2	9907	1	5873			
2	9908	1	5873			
2	9909	1	5873			
2	9910	1	5879			
2	9911	1	5879			
2	9912	1	5882			
2	9913	1	5882			
2	9914	1	5882			
2	9915	1	5886			
2	9916	1	5886			
2	9917	1	5886			
2	9918	1	5892			
2	9919	1	5892			
2	9920	1	5895			
2	9921	1	5895			
2	9922	1	5898			
2	9923	1	5898			
2	9924	1	5898			
2	9925	1	5904			
2	9926	1	5904			
2	9927	1	5907			
2	9928	1	5907			
2	9929	1	5907			
2	9930	1	5913			
2	9931	1	5913			
2	9932	1	5916			
2	9933	1	5916			
2	9934	1	5919			
2	9935	1	5919			
2	9936	1	5919			
2	9937	1	5925			
2	9938	1	5925			
2	9939	1	5930			
2	9940	1	5930			
2	9941	1	5935			
2	9942	1	5935			
2	9943	1	5938			
2	9944	1	5938			
2	9945	1	5941			
2	9946	1	5941			
2	9947	1	5941			
2	9948	1	5947			
2	9949	1	5947			
2	9950	1	5950			
2	9951	1	5950			
2	9952	1	5950			
2	9953	1	5956			
2	9954	1	5956			
2	9955	1	5959			
2	9956	1	5959			
2	9957	1	5962			
2	9958	1	5962			
2	9959	1	5962			
2	9960	1	5968			
2	9961	1	5968			
2	9962	1	5972			
2	9963	1	5972			
2	9964	1	5975			
2	9965	1	5975			
2	9966	1	5975			
2	9967	1	5981			
2	9968	1	5981			
2	9969	1	5984			
2	9970	1	5984			
2	9971	1	5984			
2	9972	1	5990			
2	9973	1	5990			
2	9974	1	5993			
2	9975	1	5993			
2	9976	1	5996			
2	9977	1	5996			
2	9978	1	5996			
2	9979	1	6002			
2	9980	1	6002			
2	9981	1	6005			
2	9982	1	6005			
2	9983	1	6005			
2	9984	1	6011			
2	9985	1	6011			
2	9986	1	6014			
2	9987	1	6014			
2	9988	1	6014			
2	9989	1	6020			
2	9990	1	6020			
2	9991	1	6023			
2	9992	1	6023			
2	9993	1	6026			
2	9994	1	6026			
2	9995	1	6026			
2	9996	1	6032			
2	9997	1	6032			
2	9998	1	6037			
2	9999	1	6037			
2	10000	1	6040			
2	10001	1	6040			
2	10002	1	6040			
2	10003	1	6046			
2	10004	1	6046			
2	10005	1	6049			
2	10006	1	6049			
2	10007	1	6052			
2	10008	1	6052			
2	10009	1	6052			
2	10010	1	6058			
2	10011	1	6058			
2	10012	1	6061			
2	10013	1	6061			
2	10014	1	6064			
2	10015	1	6064			
2	10016	1	6064			
2	10017	1	6070			
2	10018	1	6070			
2	10019	1	6073			
2	10020	1	6073			
2	10021	1	6076			
2	10022	1	6076			
2	10023	1	6076			
2	10024	1	6082			
2	10025	1	6082			
2	10026	1	6085			
2	10027	1	6085			
2	10028	1	6085			
2	10029	1	6091			
2	10030	1	6091			
2	10031	1	6094			
2	10032	1	6094			
2	10033	1	6097			
2	10034	1	6097			
2	10035	1	6097			
2	10036	1	6103			
2	10037	1	6103			
2	10038	1	6108			
2	10039	1	6108			
2	10040	1	6111			
2	10041	1	6111			
2	10042	1	6114			
2	10043	1	6114			
2	10044	1	6114			
2	10045	1	6120			
2	10046	1	6120			
2	10047	1	6124			
2	10048	1	6124			
2	10049	1	6124			
2	10050	1	6130			
2	10051	1	6130			
2	10052	1	6135			
2	10053	1	6135			
2	10054	1	6138			
2	10055	1	6138			
2	10056	1	6141			
2	10057	1	6141			
2	10058	1	6141			
2	10059	1	6147			
2	10060	1	6147			
2	10061	1	6151			
2	10062	1	6151			
2	10063	1	6151			
2	10064	1	6157			
2	10065	1	6157			
2	10066	1	6161			
2	10067	1	6161			
2	10068	1	6161			
2	10069	1	6167			
2	10070	1	6167			
2	10071	1	6171			
2	10072	1	6171			
2	10073	1	6171			
2	10074	1	6177			
2	10075	1	6177			
2	10076	1	6181			
2	10077	1	6181			
2	10078	1	6181			
2	10079	1	6187			
2	10080	1	6187			
2	10081	1	6191			
2	10082	1	6191			
2	10083	1	6191			
2	10084	1	6197			
2	10085	1	6197			
2	10086	1	6201			
2	10087	1	6201			
2	10088	1	6201			
2	10089	1	6207			
2	10090	1	6207			
2	10091	1	6211			
2	10092	1	6211			
2	10093	1	6211			
2	10094	1	6217			
2	10095	1	6217			
2	10096	1	6221			
2	10097	1	6221			
2	10098	1	6221			
2	10099	1	6227			
2	10100	1	6227			
2	10101	1	6231			
2	10102	1	6231			
2	10103	1	6231			
2	10104	1	6237			
2	10105	1	6237			
2	10106	1	6241			
2	10107	1	6241			
2	10108	1	6241			
2	10109	1	6247			
2	10110	1	6247			
2	10111	1	6251			
2	10112	1	6251			
2	10113	1	6251			
2	10114	1	6257			
2	10115	1	6257			
2	10116	1	6261			
2	10117	1	6261			
2	10118	1	6261			
2	10119	1	6267			
2	10120	1	6267			
2	10121	1	6271			
2	10122	1	6271			
2	10123	1	6271			
2	10124	1	6277			
2	10125	1	6277			
2	10126	1	6281			
2	10127	1	6281			
2	10128	1	6281			
