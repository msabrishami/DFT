1	1	0	2	0	
1	4	0	3	0	
1	8	0	2	0	
1	11	0	2	0	
1	14	0	2	0	
1	17	0	3	0	
1	21	0	2	0	
1	24	0	2	0	
1	27	0	2	0	
1	30	0	3	0	
1	34	0	2	0	
1	37	0	2	0	
1	40	0	2	0	
1	43	0	3	0	
1	47	0	2	0	
1	50	0	2	0	
1	53	0	2	0	
1	56	0	3	0	
1	60	0	2	0	
1	63	0	2	0	
1	66	0	2	0	
1	69	0	3	0	
1	73	0	2	0	
1	76	0	2	0	
1	79	0	2	0	
1	82	0	3	0	
1	86	0	2	0	
1	89	0	2	0	
1	92	0	2	0	
1	95	0	3	0	
1	99	0	2	0	
1	102	0	2	0	
1	105	0	2	0	
1	108	0	3	0	
1	112	0	2	0	
1	115	0	2	0	
0	118	5	1	1	433	
0	119	5	2	1	435	
0	122	5	1	1	440	
0	123	5	2	1	444	
0	126	5	1	1	449	
0	127	5	2	1	453	
0	130	5	1	1	458	
0	131	5	2	1	462	
0	134	5	1	1	467	
0	135	5	2	1	471	
0	138	5	1	1	476	
0	139	5	2	1	480	
0	142	5	1	1	485	
0	143	5	2	1	489	
0	146	5	1	1	494	
0	147	5	2	1	498	
0	150	5	1	1	503	
0	151	5	2	1	507	
0	154	6	2	2	118	436	
0	157	4	1	2	438	514	
0	158	4	1	2	442	515	
0	159	6	2	2	122	445	
0	162	6	2	2	126	454	
0	165	6	2	2	130	463	
0	168	6	2	2	134	472	
0	171	6	2	2	138	481	
0	174	6	2	2	142	490	
0	177	6	2	2	146	499	
0	180	6	2	2	150	508	
0	183	4	1	2	447	516	
0	184	4	1	2	451	517	
0	185	4	1	2	456	518	
0	186	4	1	2	460	519	
0	187	4	1	2	465	520	
0	188	4	1	2	469	521	
0	189	4	1	2	474	522	
0	190	4	1	2	478	523	
0	191	4	1	2	483	524	
0	192	4	1	2	487	525	
0	193	4	1	2	492	526	
0	194	4	1	2	496	527	
0	195	4	1	2	501	528	
0	196	4	1	2	505	529	
0	197	4	1	2	510	530	
0	198	4	1	2	512	531	
0	199	7	3	9	532	534	536	538	540	542	544	546	548	
0	203	5	9	1	550	
0	213	5	9	1	551	
3	223	5	0	1	552	
0	224	2	2	2	553	533	
0	227	2	2	2	554	535	
0	230	2	2	2	555	537	
0	233	2	2	2	556	539	
0	236	2	2	2	557	541	
0	239	2	2	2	558	543	
0	242	6	1	2	434	562	
0	243	2	2	2	559	545	
0	246	6	1	2	563	441	
0	247	2	2	2	560	547	
0	250	6	1	2	564	450	
0	251	2	2	2	561	549	
0	254	6	1	2	565	459	
0	255	6	1	2	566	468	
0	256	6	1	2	567	477	
0	257	6	1	2	568	486	
0	258	6	1	2	569	495	
0	259	6	1	2	570	504	
0	260	6	2	2	571	157	
0	263	6	1	2	572	158	
0	264	6	2	2	573	183	
0	267	6	2	2	575	185	
0	270	6	2	2	577	187	
0	273	6	2	2	579	189	
0	276	6	2	2	581	191	
0	279	6	2	2	583	193	
0	282	6	2	2	585	195	
0	285	6	2	2	587	197	
0	288	6	1	2	574	184	
0	289	6	1	2	576	186	
0	290	6	1	2	578	188	
0	291	6	1	2	580	190	
0	292	6	1	2	582	192	
0	293	6	1	2	584	194	
0	294	6	1	2	586	196	
0	295	6	1	2	588	198	
0	296	7	3	9	589	591	593	595	597	599	601	603	605	
0	300	5	1	1	263	
0	301	5	1	1	288	
0	302	5	1	1	289	
0	303	5	1	1	290	
0	304	5	1	1	291	
0	305	5	1	1	292	
0	306	5	1	1	293	
0	307	5	1	1	294	
0	308	5	1	1	295	
0	309	5	9	1	607	
0	319	5	9	1	608	
3	329	5	0	1	609	
0	330	2	1	2	610	590	
0	331	2	1	2	611	592	
0	332	2	1	2	612	594	
0	333	2	1	2	613	596	
0	334	6	1	2	439	619	
0	335	2	1	2	614	598	
0	336	6	1	2	620	448	
0	337	2	1	2	615	600	
0	338	6	1	2	621	457	
0	339	2	1	2	616	602	
0	340	6	1	2	622	466	
0	341	2	1	2	617	604	
0	342	6	1	2	623	475	
0	343	2	1	2	618	606	
0	344	6	1	2	624	484	
0	345	6	1	2	625	493	
0	346	6	1	2	626	502	
0	347	6	1	2	627	511	
0	348	6	1	2	330	300	
0	349	6	1	2	331	301	
0	350	6	1	2	332	302	
0	351	6	1	2	333	303	
0	352	6	1	2	335	304	
0	353	6	1	2	337	305	
0	354	6	1	2	339	306	
0	355	6	1	2	341	307	
0	356	6	1	2	343	308	
0	357	7	2	9	348	349	350	351	352	353	354	355	356	
0	360	5	9	1	628	
3	370	5	0	1	629	
0	371	6	1	2	443	630	
0	372	6	1	2	631	452	
0	373	6	1	2	632	461	
0	374	6	1	2	633	470	
0	375	6	1	2	634	479	
0	376	6	1	2	635	488	
0	377	6	1	2	636	497	
0	378	6	1	2	637	506	
0	379	6	1	2	638	513	
0	380	6	1	4	437	242	334	371	
0	381	6	4	4	246	336	372	446	
0	386	6	6	4	250	338	373	455	
0	393	6	5	4	254	340	374	464	
0	399	6	4	4	255	342	375	473	
0	404	6	2	4	256	344	376	482	
0	407	6	3	4	257	345	377	491	
0	411	6	2	4	258	346	378	500	
0	414	6	1	4	259	347	379	509	
0	415	5	1	1	380	
0	416	7	1	8	639	643	649	654	658	660	663	414	
0	417	5	1	1	650	
0	418	5	1	1	659	
0	419	5	1	1	661	
0	420	5	1	1	664	
3	421	4	0	2	415	416	
0	422	6	2	2	644	417	
0	425	6	2	4	645	651	418	655	
0	428	6	1	3	656	652	419	
0	429	6	1	4	646	653	662	420	
3	430	6	0	4	640	647	665	657	
3	431	6	0	4	641	648	667	428	
3	432	6	0	4	642	666	668	429	
2	433	1	1			
2	434	1	1			
2	435	1	4			
2	436	1	4			
2	437	1	4			
2	438	1	8			
2	439	1	8			
2	440	1	11			
2	441	1	11			
2	442	1	14			
2	443	1	14			
2	444	1	17			
2	445	1	17			
2	446	1	17			
2	447	1	21			
2	448	1	21			
2	449	1	24			
2	450	1	24			
2	451	1	27			
2	452	1	27			
2	453	1	30			
2	454	1	30			
2	455	1	30			
2	456	1	34			
2	457	1	34			
2	458	1	37			
2	459	1	37			
2	460	1	40			
2	461	1	40			
2	462	1	43			
2	463	1	43			
2	464	1	43			
2	465	1	47			
2	466	1	47			
2	467	1	50			
2	468	1	50			
2	469	1	53			
2	470	1	53			
2	471	1	56			
2	472	1	56			
2	473	1	56			
2	474	1	60			
2	475	1	60			
2	476	1	63			
2	477	1	63			
2	478	1	66			
2	479	1	66			
2	480	1	69			
2	481	1	69			
2	482	1	69			
2	483	1	73			
2	484	1	73			
2	485	1	76			
2	486	1	76			
2	487	1	79			
2	488	1	79			
2	489	1	82			
2	490	1	82			
2	491	1	82			
2	492	1	86			
2	493	1	86			
2	494	1	89			
2	495	1	89			
2	496	1	92			
2	497	1	92			
2	498	1	95			
2	499	1	95			
2	500	1	95			
2	501	1	99			
2	502	1	99			
2	503	1	102			
2	504	1	102			
2	505	1	105			
2	506	1	105			
2	507	1	108			
2	508	1	108			
2	509	1	108			
2	510	1	112			
2	511	1	112			
2	512	1	115			
2	513	1	115			
2	514	1	119			
2	515	1	119			
2	516	1	123			
2	517	1	123			
2	518	1	127			
2	519	1	127			
2	520	1	131			
2	521	1	131			
2	522	1	135			
2	523	1	135			
2	524	1	139			
2	525	1	139			
2	526	1	143			
2	527	1	143			
2	528	1	147			
2	529	1	147			
2	530	1	151			
2	531	1	151			
2	532	1	154			
2	533	1	154			
2	534	1	159			
2	535	1	159			
2	536	1	162			
2	537	1	162			
2	538	1	165			
2	539	1	165			
2	540	1	168			
2	541	1	168			
2	542	1	171			
2	543	1	171			
2	544	1	174			
2	545	1	174			
2	546	1	177			
2	547	1	177			
2	548	1	180			
2	549	1	180			
2	550	1	199			
2	551	1	199			
2	552	1	199			
2	553	1	203			
2	554	1	203			
2	555	1	203			
2	556	1	203			
2	557	1	203			
2	558	1	203			
2	559	1	203			
2	560	1	203			
2	561	1	203			
2	562	1	213			
2	563	1	213			
2	564	1	213			
2	565	1	213			
2	566	1	213			
2	567	1	213			
2	568	1	213			
2	569	1	213			
2	570	1	213			
2	571	1	224			
2	572	1	224			
2	573	1	227			
2	574	1	227			
2	575	1	230			
2	576	1	230			
2	577	1	233			
2	578	1	233			
2	579	1	236			
2	580	1	236			
2	581	1	239			
2	582	1	239			
2	583	1	243			
2	584	1	243			
2	585	1	247			
2	586	1	247			
2	587	1	251			
2	588	1	251			
2	589	1	260			
2	590	1	260			
2	591	1	264			
2	592	1	264			
2	593	1	267			
2	594	1	267			
2	595	1	270			
2	596	1	270			
2	597	1	273			
2	598	1	273			
2	599	1	276			
2	600	1	276			
2	601	1	279			
2	602	1	279			
2	603	1	282			
2	604	1	282			
2	605	1	285			
2	606	1	285			
2	607	1	296			
2	608	1	296			
2	609	1	296			
2	610	1	309			
2	611	1	309			
2	612	1	309			
2	613	1	309			
2	614	1	309			
2	615	1	309			
2	616	1	309			
2	617	1	309			
2	618	1	309			
2	619	1	319			
2	620	1	319			
2	621	1	319			
2	622	1	319			
2	623	1	319			
2	624	1	319			
2	625	1	319			
2	626	1	319			
2	627	1	319			
2	628	1	357			
2	629	1	357			
2	630	1	360			
2	631	1	360			
2	632	1	360			
2	633	1	360			
2	634	1	360			
2	635	1	360			
2	636	1	360			
2	637	1	360			
2	638	1	360			
2	639	1	381			
2	640	1	381			
2	641	1	381			
2	642	1	381			
2	643	1	386			
2	644	1	386			
2	645	1	386			
2	646	1	386			
2	647	1	386			
2	648	1	386			
2	649	1	393			
2	650	1	393			
2	651	1	393			
2	652	1	393			
2	653	1	393			
2	654	1	399			
2	655	1	399			
2	656	1	399			
2	657	1	399			
2	658	1	404			
2	659	1	404			
2	660	1	407			
2	661	1	407			
2	662	1	407			
2	663	1	411			
2	664	1	411			
2	665	1	422			
2	666	1	422			
2	667	1	425			
2	668	1	425			
