<<<<<<< HEAD
1 1 0 2 0
2 13 1 1
2 14 1 1
1 4 0 3 0
2 15 1 4
2 16 1 4
2 17 1 4
1 8 0 3 0
2 18 1 8
2 19 1 8
2 20 1 8
1 12 0 2 0
2 21 1 12
2 22 1 12
0 23 6 1 2 13 18
0 24 6 2 2 16 19
2 28 1 24 
2 29 1 24
0 27 6 1 2 17 22
0 30 6 1 2 15 23
0 31 6 1 2 14 28
0 32 6 1 2 29 21
0 33 6 1 2 27 20
=======
1 1 0 2 0
2 13 1 1
2 14 1 1
1 4 0 3 0
2 15 1 4
2 16 1 4
2 17 1 4
1 8 0 3 0
2 18 1 8
2 19 1 8
2 20 1 8
1 12 0 2 0
2 21 1 12
2 22 1 12
0 23 6 1 2 13 18
0 24 6 2 2 16 19
2 28 1 24 
2 29 1 24
0 27 6 1 2 17 22
0 30 6 1 2 15 23
0 31 6 1 2 14 28
0 32 6 1 2 29 21
0 33 6 1 2 27 20
>>>>>>> 8b13aad36fc8e5900215a2790ecd424518d66181
3 34 6 0 4 30 31 32 33