1	1	0	6	0	
1	8	0	4	0	
1	13	0	3	0	
1	17	0	8	0	
1	26	0	2	0	
1	29	0	6	0	
1	36	0	5	0	
1	42	0	8	0	
1	51	0	3	0	
1	55	0	3	0	
1	59	0	8	0	
1	68	0	3	0	
1	72	0	1	0	
1	73	0	1	0	
1	74	0	1	0	
1	75	0	4	0	
1	80	0	4	0	
1	85	0	1	0	
1	86	0	1	0	
1	87	0	1	0	
1	88	0	1	0	
1	89	0	1	0	
1	90	0	1	0	
1	91	0	4	0	
1	96	0	4	0	
1	101	0	4	0	
1	106	0	4	0	
1	111	0	4	0	
1	116	0	4	0	
1	121	0	4	0	
1	126	0	3	0	
1	130	0	4	0	
1	135	0	2	0	
1	138	0	4	0	
1	143	0	2	0	
1	146	0	2	0	
1	149	0	2	0	
1	152	0	1	0	
1	153	0	2	0	
1	156	0	2	0	
1	159	0	5	0	
1	165	0	5	0	
1	171	0	5	0	
1	177	0	5	0	
1	183	0	5	0	
1	189	0	5	0	
1	195	0	5	0	
1	201	0	5	0	
1	207	0	2	0	
1	210	0	8	0	
1	219	0	8	0	
1	228	0	8	0	
1	237	0	8	0	
1	246	0	8	0	
1	255	0	3	0	
1	259	0	1	0	
1	260	0	1	0	
1	261	0	5	0	
1	267	0	1	0	
1	268	0	1	0	
0	269	6	1	4	878	884	888	891	
0	270	6	2	4	879	899	889	892	
0	273	7	2	3	901	907	912	
0	276	7	2	3	880	900	920	
0	279	6	1	4	881	885	921	893	
0	280	6	3	4	882	886	890	923	
0	284	6	1	4	926	913	934	72	
0	285	6	1	2	902	935	
0	286	6	1	3	927	936	74	
0	287	7	2	3	903	937	941	
3	290	7	0	3	904	938	914	
3	291	7	0	3	905	908	942	
3	292	7	0	3	906	909	915	
0	293	7	1	3	928	939	943	
0	294	7	1	3	929	940	916	
0	295	7	1	3	930	910	944	
0	296	7	1	3	931	911	917	
3	297	7	0	2	85	86	
0	298	3	2	2	87	88	
0	301	6	1	2	945	949	
0	302	3	1	2	946	950	
0	303	6	1	2	953	957	
0	304	3	1	2	954	958	
0	305	6	1	2	961	965	
0	306	3	1	2	962	966	
0	307	6	1	2	969	973	
0	308	3	1	2	970	974	
0	309	7	1	2	887	982	
0	310	5	5	1	268	
0	316	7	1	2	922	983	
0	317	7	1	2	894	984	
0	318	7	1	2	152	985	
0	319	6	2	2	932	994	
0	322	4	1	2	895	918	
0	323	7	1	2	896	919	
0	324	6	1	2	996	1001	
0	325	3	1	2	997	1002	
0	326	6	1	2	1006	1011	
0	327	3	1	2	1007	1012	
0	328	6	1	2	1016	1021	
0	329	3	1	2	1017	1022	
0	330	6	1	2	1026	1031	
0	331	3	1	2	1027	1032	
0	332	7	1	2	1038	947	
0	333	7	1	2	1039	951	
0	334	7	1	2	1040	955	
0	335	7	1	2	1041	959	
0	336	7	1	2	1042	963	
0	337	7	1	2	1078	259	
0	338	7	1	2	1043	967	
0	339	7	1	2	1079	260	
0	340	7	1	2	1044	971	
0	341	7	1	2	1080	267	
3	342	5	0	1	269	
0	343	5	1	1	1088	
3	344	3	0	2	1086	1089	
0	345	5	1	1	1090	
0	346	5	1	1	1091	
0	347	5	1	1	279	
0	348	4	1	2	1092	284	
0	349	3	1	2	1093	285	
0	350	3	1	2	1094	286	
3	351	5	0	1	293	
0	352	5	1	1	294	
3	353	5	0	1	295	
3	354	5	0	1	296	
0	355	6	1	2	89	1097	
3	356	7	0	2	90	1098	
0	357	6	2	2	301	302	
0	360	6	2	2	303	304	
0	363	6	2	2	305	306	
0	366	6	2	2	307	308	
0	369	5	5	1	1099	
0	375	4	1	2	322	323	
0	376	6	2	2	324	325	
0	379	6	2	2	326	327	
0	382	6	2	2	328	329	
0	385	6	2	2	330	331	
3	392	3	0	2	1087	343	
0	393	5	5	1	345	
3	399	5	0	1	346	
0	400	7	1	2	348	73	
3	401	5	0	1	349	
3	402	5	0	1	350	
3	403	5	0	1	355	
0	404	5	1	1	1106	
0	405	5	1	1	1108	
0	406	7	1	2	1107	1109	
0	407	5	1	1	1110	
0	408	5	1	1	1112	
0	409	7	1	2	1111	1113	
0	410	6	1	2	347	352	
0	411	5	1	1	1119	
0	412	5	1	1	1121	
0	413	7	1	2	1120	1122	
0	414	5	1	1	1123	
0	415	5	1	1	1125	
0	416	7	1	2	1124	1126	
0	417	7	1	2	1045	1114	
0	424	5	1	1	400	
0	425	7	1	2	404	405	
0	426	7	1	2	407	408	
0	427	7	4	3	1104	1127	924	
0	432	7	4	3	1128	897	1095	
0	437	6	4	3	1129	1096	925	
0	442	6	1	4	375	933	995	1130	
0	443	6	1	3	1131	1105	898	
0	444	7	1	2	411	412	
0	445	7	1	2	414	415	
0	451	5	8	1	424	
0	460	4	2	2	406	425	
0	463	4	2	2	409	426	
0	466	6	8	2	442	410	
0	475	7	1	2	986	1132	
0	476	7	1	2	1100	1136	
0	477	7	1	2	988	1133	
0	478	7	1	2	1101	1137	
0	479	7	1	2	990	1134	
0	480	7	1	2	1102	1138	
0	481	7	1	2	992	1135	
0	482	7	1	2	1103	1139	
0	483	6	4	2	443	883	
0	488	3	1	2	1115	1140	
0	489	3	1	2	1116	1141	
0	490	3	1	2	1117	1142	
0	491	3	1	2	1118	1143	
0	492	4	2	2	413	444	
0	495	4	2	2	416	445	
0	498	6	1	2	976	1152	
0	499	3	1	2	977	1153	
0	500	6	1	2	1154	980	
0	501	3	1	2	1155	981	
0	502	7	1	2	948	1156	
0	503	4	1	2	475	476	
0	504	7	1	2	952	1157	
0	505	4	1	2	477	478	
0	506	7	1	2	956	1158	
0	507	4	1	2	479	480	
0	508	7	1	2	960	1159	
0	509	4	1	2	481	482	
0	510	7	1	2	987	1164	
0	511	7	1	2	964	1160	
0	512	7	1	2	989	1165	
0	513	7	1	2	968	1161	
0	514	7	1	2	991	1166	
0	515	7	1	2	972	1162	
0	516	7	1	2	993	1167	
0	517	7	1	2	975	1163	
0	518	6	1	2	978	1168	
0	519	3	1	2	979	1169	
0	520	6	1	2	1170	1036	
0	521	3	1	2	1171	1037	
0	522	7	1	2	1144	998	
0	523	7	1	2	1145	1003	
0	524	7	1	2	1146	1008	
0	525	7	1	2	1147	1013	
0	526	7	1	2	1148	1018	
0	527	6	1	2	1149	1023	
0	528	6	1	2	1150	1028	
0	529	6	1	2	1151	1033	
0	530	6	2	2	498	499	
0	533	6	2	2	500	501	
0	536	4	1	2	309	502	
0	537	4	1	2	316	504	
0	538	4	1	2	317	506	
0	539	4	1	2	318	508	
0	540	4	1	2	510	511	
0	541	4	1	2	512	513	
0	542	4	1	2	514	515	
0	543	4	1	2	516	517	
0	544	6	2	2	518	519	
0	547	6	2	2	520	521	
0	550	5	1	1	1172	
0	551	5	1	1	1174	
0	552	7	1	2	1173	1175	
0	553	6	3	2	536	503	
0	557	6	3	2	537	505	
0	561	6	3	2	538	507	
0	565	6	3	2	539	509	
0	569	6	3	2	488	540	
0	573	6	3	2	489	541	
0	577	6	3	2	490	542	
0	581	6	3	2	491	543	
0	585	5	1	1	1176	
0	586	5	1	1	1178	
0	587	7	1	2	1177	1179	
0	588	7	1	2	550	551	
0	589	7	1	2	585	586	
0	590	6	2	2	1180	999	
0	593	3	2	2	1181	1000	
0	596	7	1	2	1070	1182	
0	597	6	2	2	1183	1004	
0	600	3	4	2	1184	1005	
0	605	7	1	2	1071	1185	
0	606	6	2	2	1186	1009	
0	609	3	5	2	1187	1010	
0	615	7	1	2	1072	1188	
0	616	6	2	2	1189	1014	
0	619	3	4	2	1190	1015	
0	624	7	1	2	1073	1191	
0	625	6	2	2	1192	1019	
0	628	3	2	2	1193	1020	
0	631	7	1	2	1074	1194	
0	632	6	2	2	1195	1024	
0	635	3	4	2	1196	1025	
0	640	7	1	2	1075	1197	
0	641	6	2	2	1198	1029	
0	644	3	5	2	1199	1030	
0	650	7	1	2	1076	1200	
0	651	6	2	2	1201	1034	
0	654	3	4	2	1202	1035	
0	659	7	1	2	1077	1203	
3	660	4	0	2	552	588	
3	661	4	0	2	587	589	
0	662	5	2	1	1204	
0	665	7	3	2	1206	1205	
0	669	4	1	2	596	522	
0	670	5	2	1	1208	
0	673	7	3	2	1210	1209	
0	677	4	1	2	605	523	
0	678	5	3	1	1214	
0	682	7	3	2	1216	1215	
0	686	4	1	2	615	524	
0	687	5	4	1	1221	
0	692	7	3	2	1223	1222	
0	696	4	1	2	624	525	
0	697	5	2	1	1227	
0	700	7	3	2	1229	1228	
0	704	4	1	2	631	526	
0	705	5	2	1	1231	
0	708	7	3	2	1233	1232	
0	712	4	1	2	337	640	
0	713	5	3	1	1237	
0	717	7	3	2	1239	1238	
0	721	4	1	2	339	650	
0	722	5	4	1	1244	
0	727	7	3	2	1246	1245	
0	731	4	1	2	341	659	
0	732	6	1	2	1247	1081	
0	733	6	1	3	1240	1248	1082	
0	734	6	1	4	1234	1241	1249	1083	
0	735	5	1	1	1250	
0	736	7	1	2	1054	1252	
0	737	7	1	2	1062	1251	
0	738	5	1	1	1255	
0	739	7	1	2	1055	1257	
0	740	7	1	2	1063	1256	
0	741	5	1	1	1260	
0	742	7	1	2	1056	1263	
0	743	7	1	2	1064	1261	
0	744	5	1	1	1266	
0	745	7	1	2	1057	1270	
0	746	7	1	2	1065	1267	
0	747	5	1	1	1273	
0	748	7	1	2	1058	1275	
0	749	7	1	2	1066	1274	
0	750	5	1	1	1278	
0	751	7	1	2	1059	1280	
0	752	7	1	2	1067	1279	
0	753	5	1	1	1283	
0	754	7	1	2	1060	1286	
0	755	7	1	2	1068	1284	
0	756	5	1	1	1289	
0	757	4	1	2	1293	1084	
0	758	7	1	2	1294	1085	
0	759	7	1	2	1061	1295	
0	760	7	1	2	1069	1290	
0	761	6	1	2	1242	1291	
0	762	6	1	2	1235	1285	
0	763	6	1	3	1236	1243	1292	
0	764	6	1	2	1217	1268	
0	765	6	1	2	1211	1262	
0	766	6	1	3	1212	1218	1269	
0	769	4	1	2	736	737	
0	770	4	1	2	739	740	
0	771	4	1	2	742	743	
0	772	4	1	2	745	746	
0	773	6	3	4	750	762	763	734	
0	777	4	1	2	748	749	
0	778	6	2	3	753	761	733	
0	781	4	1	2	751	752	
0	782	6	2	2	756	732	
0	785	4	1	2	754	755	
0	786	4	1	2	757	758	
0	787	4	1	2	759	760	
0	788	4	1	2	1276	1296	
0	789	7	1	2	1277	1297	
0	790	4	1	2	1281	1299	
0	791	7	1	2	1282	1300	
0	792	4	1	2	1287	1301	
0	793	7	1	2	1288	1302	
0	794	7	1	2	1046	786	
0	795	6	1	2	1230	1298	
0	796	6	5	2	795	747	
0	802	4	1	2	788	789	
0	803	4	1	2	790	791	
0	804	4	1	2	792	793	
0	805	4	1	2	340	794	
0	806	4	1	2	1271	1303	
0	807	7	1	2	1272	1304	
0	808	7	1	2	1047	802	
0	809	7	1	2	1048	803	
0	810	7	1	2	1049	804	
0	811	6	1	4	805	787	731	529	
0	812	6	1	2	1224	1305	
0	813	6	1	3	1219	1225	1306	
0	814	6	1	4	1213	1220	1226	1307	
0	815	6	3	4	738	765	766	814	
0	819	6	2	3	741	764	813	
0	822	6	2	2	744	812	
0	825	4	1	2	806	807	
0	826	4	1	2	335	808	
0	827	4	1	2	336	809	
0	828	4	1	2	338	810	
0	829	5	1	1	811	
0	830	4	1	2	1253	1308	
0	831	7	1	2	1254	1309	
0	832	4	1	2	1258	1311	
0	833	7	1	2	1259	1312	
0	834	4	1	2	1264	1313	
0	835	7	1	2	1265	1314	
0	836	7	1	2	1050	825	
0	837	6	1	3	826	777	704	
0	838	6	1	4	827	781	712	527	
0	839	6	1	4	828	785	721	528	
3	840	5	0	1	829	
0	841	6	1	2	1310	1207	
0	842	4	1	2	830	831	
0	843	4	1	2	832	833	
0	844	4	1	2	834	835	
0	845	4	1	2	334	836	
0	846	5	1	1	837	
0	847	5	1	1	838	
0	848	5	1	1	839	
0	849	7	1	2	735	841	
0	851	7	1	2	1051	842	
0	852	7	1	2	1052	843	
0	853	7	1	2	1053	844	
0	854	6	1	3	845	772	696	
3	855	5	0	1	846	
3	856	5	0	1	847	
3	857	5	0	1	848	
3	858	5	0	1	849	
0	859	4	1	2	417	851	
0	860	4	1	2	332	852	
0	861	4	1	2	333	853	
0	862	5	1	1	854	
0	867	6	1	3	859	769	669	
0	868	6	1	3	860	770	677	
0	869	6	1	3	861	771	686	
3	870	5	0	1	862	
0	871	5	1	1	867	
0	872	5	1	1	868	
0	873	5	1	1	869	
3	875	5	0	1	871	
3	876	5	0	1	872	
3	877	5	0	1	873	
2	878	1	1			
2	879	1	1			
2	880	1	1			
2	881	1	1			
2	882	1	1			
2	883	1	1			
2	884	1	8			
2	885	1	8			
2	886	1	8			
2	887	1	8			
2	888	1	13			
2	889	1	13			
2	890	1	13			
2	891	1	17			
2	892	1	17			
2	893	1	17			
2	894	1	17			
2	895	1	17			
2	896	1	17			
2	897	1	17			
2	898	1	17			
2	899	1	26			
2	900	1	26			
2	901	1	29			
2	902	1	29			
2	903	1	29			
2	904	1	29			
2	905	1	29			
2	906	1	29			
2	907	1	36			
2	908	1	36			
2	909	1	36			
2	910	1	36			
2	911	1	36			
2	912	1	42			
2	913	1	42			
2	914	1	42			
2	915	1	42			
2	916	1	42			
2	917	1	42			
2	918	1	42			
2	919	1	42			
2	920	1	51			
2	921	1	51			
2	922	1	51			
2	923	1	55			
2	924	1	55			
2	925	1	55			
2	926	1	59			
2	927	1	59			
2	928	1	59			
2	929	1	59			
2	930	1	59			
2	931	1	59			
2	932	1	59			
2	933	1	59			
2	934	1	68			
2	935	1	68			
2	936	1	68			
2	937	1	75			
2	938	1	75			
2	939	1	75			
2	940	1	75			
2	941	1	80			
2	942	1	80			
2	943	1	80			
2	944	1	80			
2	945	1	91			
2	946	1	91			
2	947	1	91			
2	948	1	91			
2	949	1	96			
2	950	1	96			
2	951	1	96			
2	952	1	96			
2	953	1	101			
2	954	1	101			
2	955	1	101			
2	956	1	101			
2	957	1	106			
2	958	1	106			
2	959	1	106			
2	960	1	106			
2	961	1	111			
2	962	1	111			
2	963	1	111			
2	964	1	111			
2	965	1	116			
2	966	1	116			
2	967	1	116			
2	968	1	116			
2	969	1	121			
2	970	1	121			
2	971	1	121			
2	972	1	121			
2	973	1	126			
2	974	1	126			
2	975	1	126			
2	976	1	130			
2	977	1	130			
2	978	1	130			
2	979	1	130			
2	980	1	135			
2	981	1	135			
2	982	1	138			
2	983	1	138			
2	984	1	138			
2	985	1	138			
2	986	1	143			
2	987	1	143			
2	988	1	146			
2	989	1	146			
2	990	1	149			
2	991	1	149			
2	992	1	153			
2	993	1	153			
2	994	1	156			
2	995	1	156			
2	996	1	159			
2	997	1	159			
2	998	1	159			
2	999	1	159			
2	1000	1	159			
2	1001	1	165			
2	1002	1	165			
2	1003	1	165			
2	1004	1	165			
2	1005	1	165			
2	1006	1	171			
2	1007	1	171			
2	1008	1	171			
2	1009	1	171			
2	1010	1	171			
2	1011	1	177			
2	1012	1	177			
2	1013	1	177			
2	1014	1	177			
2	1015	1	177			
2	1016	1	183			
2	1017	1	183			
2	1018	1	183			
2	1019	1	183			
2	1020	1	183			
2	1021	1	189			
2	1022	1	189			
2	1023	1	189			
2	1024	1	189			
2	1025	1	189			
2	1026	1	195			
2	1027	1	195			
2	1028	1	195			
2	1029	1	195			
2	1030	1	195			
2	1031	1	201			
2	1032	1	201			
2	1033	1	201			
2	1034	1	201			
2	1035	1	201			
2	1036	1	207			
2	1037	1	207			
2	1038	1	210			
2	1039	1	210			
2	1040	1	210			
2	1041	1	210			
2	1042	1	210			
2	1043	1	210			
2	1044	1	210			
2	1045	1	210			
2	1046	1	219			
2	1047	1	219			
2	1048	1	219			
2	1049	1	219			
2	1050	1	219			
2	1051	1	219			
2	1052	1	219			
2	1053	1	219			
2	1054	1	228			
2	1055	1	228			
2	1056	1	228			
2	1057	1	228			
2	1058	1	228			
2	1059	1	228			
2	1060	1	228			
2	1061	1	228			
2	1062	1	237			
2	1063	1	237			
2	1064	1	237			
2	1065	1	237			
2	1066	1	237			
2	1067	1	237			
2	1068	1	237			
2	1069	1	237			
2	1070	1	246			
2	1071	1	246			
2	1072	1	246			
2	1073	1	246			
2	1074	1	246			
2	1075	1	246			
2	1076	1	246			
2	1077	1	246			
2	1078	1	255			
2	1079	1	255			
2	1080	1	255			
2	1081	1	261			
2	1082	1	261			
2	1083	1	261			
2	1084	1	261			
2	1085	1	261			
2	1086	1	270			
2	1087	1	270			
2	1088	1	273			
2	1089	1	273			
2	1090	1	276			
2	1091	1	276			
2	1092	1	280			
2	1093	1	280			
2	1094	1	280			
2	1095	1	287			
2	1096	1	287			
2	1097	1	298			
2	1098	1	298			
2	1099	1	310			
2	1100	1	310			
2	1101	1	310			
2	1102	1	310			
2	1103	1	310			
2	1104	1	319			
2	1105	1	319			
2	1106	1	357			
2	1107	1	357			
2	1108	1	360			
2	1109	1	360			
2	1110	1	363			
2	1111	1	363			
2	1112	1	366			
2	1113	1	366			
2	1114	1	369			
2	1115	1	369			
2	1116	1	369			
2	1117	1	369			
2	1118	1	369			
2	1119	1	376			
2	1120	1	376			
2	1121	1	379			
2	1122	1	379			
2	1123	1	382			
2	1124	1	382			
2	1125	1	385			
2	1126	1	385			
2	1127	1	393			
2	1128	1	393			
2	1129	1	393			
2	1130	1	393			
2	1131	1	393			
2	1132	1	427			
2	1133	1	427			
2	1134	1	427			
2	1135	1	427			
2	1136	1	432			
2	1137	1	432			
2	1138	1	432			
2	1139	1	432			
2	1140	1	437			
2	1141	1	437			
2	1142	1	437			
2	1143	1	437			
2	1144	1	451			
2	1145	1	451			
2	1146	1	451			
2	1147	1	451			
2	1148	1	451			
2	1149	1	451			
2	1150	1	451			
2	1151	1	451			
2	1152	1	460			
2	1153	1	460			
2	1154	1	463			
2	1155	1	463			
2	1156	1	466			
2	1157	1	466			
2	1158	1	466			
2	1159	1	466			
2	1160	1	466			
2	1161	1	466			
2	1162	1	466			
2	1163	1	466			
2	1164	1	483			
2	1165	1	483			
2	1166	1	483			
2	1167	1	483			
2	1168	1	492			
2	1169	1	492			
2	1170	1	495			
2	1171	1	495			
2	1172	1	530			
2	1173	1	530			
2	1174	1	533			
2	1175	1	533			
2	1176	1	544			
2	1177	1	544			
2	1178	1	547			
2	1179	1	547			
2	1180	1	553			
2	1181	1	553			
2	1182	1	553			
2	1183	1	557			
2	1184	1	557			
2	1185	1	557			
2	1186	1	561			
2	1187	1	561			
2	1188	1	561			
2	1189	1	565			
2	1190	1	565			
2	1191	1	565			
2	1192	1	569			
2	1193	1	569			
2	1194	1	569			
2	1195	1	573			
2	1196	1	573			
2	1197	1	573			
2	1198	1	577			
2	1199	1	577			
2	1200	1	577			
2	1201	1	581			
2	1202	1	581			
2	1203	1	581			
2	1204	1	590			
2	1205	1	590			
2	1206	1	593			
2	1207	1	593			
2	1208	1	597			
2	1209	1	597			
2	1210	1	600			
2	1211	1	600			
2	1212	1	600			
2	1213	1	600			
2	1214	1	606			
2	1215	1	606			
2	1216	1	609			
2	1217	1	609			
2	1218	1	609			
2	1219	1	609			
2	1220	1	609			
2	1221	1	616			
2	1222	1	616			
2	1223	1	619			
2	1224	1	619			
2	1225	1	619			
2	1226	1	619			
2	1227	1	625			
2	1228	1	625			
2	1229	1	628			
2	1230	1	628			
2	1231	1	632			
2	1232	1	632			
2	1233	1	635			
2	1234	1	635			
2	1235	1	635			
2	1236	1	635			
2	1237	1	641			
2	1238	1	641			
2	1239	1	644			
2	1240	1	644			
2	1241	1	644			
2	1242	1	644			
2	1243	1	644			
2	1244	1	651			
2	1245	1	651			
2	1246	1	654			
2	1247	1	654			
2	1248	1	654			
2	1249	1	654			
2	1250	1	662			
2	1251	1	662			
2	1252	1	665			
2	1253	1	665			
2	1254	1	665			
2	1255	1	670			
2	1256	1	670			
2	1257	1	673			
2	1258	1	673			
2	1259	1	673			
2	1260	1	678			
2	1261	1	678			
2	1262	1	678			
2	1263	1	682			
2	1264	1	682			
2	1265	1	682			
2	1266	1	687			
2	1267	1	687			
2	1268	1	687			
2	1269	1	687			
2	1270	1	692			
2	1271	1	692			
2	1272	1	692			
2	1273	1	697			
2	1274	1	697			
2	1275	1	700			
2	1276	1	700			
2	1277	1	700			
2	1278	1	705			
2	1279	1	705			
2	1280	1	708			
2	1281	1	708			
2	1282	1	708			
2	1283	1	713			
2	1284	1	713			
2	1285	1	713			
2	1286	1	717			
2	1287	1	717			
2	1288	1	717			
2	1289	1	722			
2	1290	1	722			
2	1291	1	722			
2	1292	1	722			
2	1293	1	727			
2	1294	1	727			
2	1295	1	727			
2	1296	1	773			
2	1297	1	773			
2	1298	1	773			
2	1299	1	778			
2	1300	1	778			
2	1301	1	782			
2	1302	1	782			
2	1303	1	796			
2	1304	1	796			
2	1305	1	796			
2	1306	1	796			
2	1307	1	796			
2	1308	1	815			
2	1309	1	815			
2	1310	1	815			
2	1311	1	819			
2	1312	1	819			
2	1313	1	822			
2	1314	1	822			
