1 0 0 2 0
1 1 0 3 0
1 2 0 3 0
1 3 0 2 0
1 4 0 2 0
1 5 0 3 0
1 6 0 1 0
1 7 0 1 0
1 8 0 2 0
1 9 0 2 0
1 10 0 2 0
1 11 0 2 0
1 12 0 2 0
1 13 0 2 0
1 14 0 2 0
1 15 0 2 0
1 16 0 2 0
1 17 0 2 0
1 18 0 1 0
1 19 0 2 0
1 20 0 2 0
1 21 0 2 0
1 22 0 1 0
1 23 0 2 0
1 24 0 2 0
1 25 0 2 0
1 26 0 2 0
1 27 0 2 0
1 28 0 1 0
1 29 0 2 0
1 30 0 1 0
1 31 0 2 0
1 32 0 1 0
1 33 0 3 0
1 34 0 1 0
1 35 0 1 0
0 36 5 2 1 28
0 37 5 2 1 32
0 38 5 2 1 30
0 39 5 2 1 6
0 40 5 2 1 22
0 41 5 2 1 18
2 42 1 0 
2 43 1 0 
2 44 1 1 
2 45 1 1 
2 46 1 1 
2 47 1 2 
2 48 1 2 
2 49 1 2 
2 50 1 3 
2 51 1 3 
2 52 1 4 
2 53 1 4 
2 54 1 5 
2 55 1 5 
2 56 1 5 
2 57 1 8 
2 58 1 8 
2 59 1 9 
2 60 1 9 
2 61 1 10 
2 62 1 10 
2 63 1 11 
2 64 1 11 
2 65 1 12 
2 66 1 12 
2 67 1 13 
2 68 1 13 
2 69 1 14 
2 70 1 14 
2 71 1 15 
2 72 1 15 
2 73 1 16 
2 74 1 16 
2 75 1 17 
2 76 1 17 
2 77 1 19 
2 78 1 19 
2 79 1 20 
2 80 1 20 
2 81 1 21 
2 82 1 21 
2 83 1 23 
2 84 1 23 
2 85 1 24 
2 86 1 24 
2 87 1 25 
2 88 1 25 
2 89 1 26 
2 90 1 26 
2 91 1 27 
2 92 1 27 
2 93 1 29 
2 94 1 29 
2 95 1 31 
2 96 1 31 
2 97 1 33 
2 98 1 33 
2 99 1 33 
0 100 5 1 1 73
0 101 5 1 1 54
0 102 5 2 1 51
0 103 5 1 1 64
0 104 5 1 1 96
0 105 5 2 1 46
0 106 5 3 1 60
0 107 5 1 1 84
0 108 5 1 1 92
0 109 5 1 1 72
0 110 5 1 1 78
2 111 1 36 
2 112 1 36 
2 113 1 37 
2 114 1 37 
2 115 1 38 
2 116 1 38 
2 117 1 39 
2 118 1 39 
2 119 1 40 
2 120 1 40 
2 121 1 41 
2 122 1 41 
0 123 6 1 2 103 68
0 124 6 1 2 104 99
0 125 6 1 2 107 88
0 126 6 1 2 108 94
0 127 6 1 2 109 76
0 128 6 1 2 110 82
2 129 1 102 
2 130 1 102 
2 131 1 105 
2 132 1 105 
2 133 1 106 
2 134 1 106 
2 135 1 106 
0 136 6 1 2 56 130
0 137 4 1 2 43 132
0 138 4 2 2 7 135
0 139 6 1 2 126 125
0 140 6 1 2 128 127
0 141 6 1 2 123 136
0 142 4 1 2 140 139
2 143 1 138 
2 144 1 138 
0 145 4 1 2 137 144
0 146 6 1 2 145 124
0 147 4 1 2 146 141
3 148 6 0 2 142 147
2 149 1 148 
2 150 1 148 
2 151 1 148 
2 152 1 148 
2 153 1 148 
2 154 1 148 
2 155 1 148 
2 156 1 148 
2 157 1 148 
0 158 6 1 2 91 149
0 159 6 1 2 50 150
0 160 6 1 2 95 151
0 161 6 1 2 77 152
0 162 6 1 2 83 153
0 163 6 1 2 63 154
0 164 6 2 2 42 155
0 165 5 2 1 156
0 166 6 1 2 71 157
0 167 6 2 2 158 93
0 168 7 2 2 159 55
0 169 6 2 2 160 98
0 170 7 3 2 161 81
0 171 6 3 2 162 87
0 172 6 3 2 163 67
0 173 7 3 2 166 75
2 174 1 164 
2 175 1 164 
2 176 1 165 
2 177 1 165 
0 178 4 1 2 176 129
0 179 5 2 1 175
0 180 4 3 2 177 143
2 181 1 167 
2 182 1 167 
2 183 1 168 
2 184 1 168 
2 185 1 169 
2 186 1 169 
2 187 1 170 
2 188 1 170 
2 189 1 170 
2 190 1 171 
2 191 1 171 
2 192 1 171 
2 193 1 172 
2 194 1 172 
2 195 1 172 
2 196 1 173 
2 197 1 173 
2 198 1 173 
0 199 5 1 1 185
0 200 5 2 1 194
0 201 4 1 2 178 101
0 202 5 2 1 182
0 203 6 2 2 118 184
0 204 4 2 2 34 186
0 205 7 2 2 120 189
0 206 4 2 2 90 192
0 207 4 3 2 70 195
0 208 6 2 2 122 198
2 209 1 179 
2 210 1 179 
2 211 1 180 
2 212 1 180 
2 213 1 180 
0 214 4 1 2 53 209
0 215 4 1 2 66 212
0 216 4 1 2 49 210
0 217 4 1 2 62 213
2 218 1 200 
2 219 1 200 
2 220 1 202 
2 221 1 202 
2 222 1 203 
2 223 1 203 
2 224 1 204 
2 225 1 204 
2 226 1 205 
2 227 1 205 
2 228 1 206 
2 229 1 206 
2 230 1 207 
2 231 1 207 
2 232 1 207 
2 233 1 208 
2 234 1 208 
0 235 6 2 2 116 221
0 236 5 1 1 225
0 237 4 1 2 227 229
0 238 5 1 1 232
0 239 6 1 2 216 45
0 240 6 2 2 217 59
0 241 6 1 2 237 236
0 242 6 1 2 239 238
2 243 1 235 
2 244 1 235 
2 245 1 240 
2 246 1 240 
0 247 6 1 2 244 223
0 248 6 1 2 246 234
0 249 4 1 2 241 247
0 250 4 1 2 248 242
3 251 6 0 2 250 249
2 252 1 251 
2 253 1 251 
2 254 1 251 
2 255 1 251 
2 256 1 251 
2 257 1 251 
2 258 1 251 
2 259 1 251 
2 260 1 251 
2 261 1 251 
2 262 1 251 
0 263 4 1 2 252 193
0 264 7 1 2 89 253
0 265 7 1 2 69 254
0 266 7 1 2 61 255
0 267 6 1 2 47 256
0 268 7 1 2 48 257
0 269 6 1 2 258 243
0 270 7 1 2 259 222
0 271 7 1 2 260 245
0 272 5 8 1 261
0 273 7 1 2 262 233
0 274 4 1 2 263 230
0 275 4 1 2 266 211
0 276 6 1 2 267 174
0 277 4 1 2 268 131
0 278 6 1 2 269 114
0 279 4 1 2 270 58
0 280 4 1 2 271 134
0 281 4 1 2 273 80
2 282 1 272 
2 283 1 272 
2 284 1 272 
2 285 1 272 
2 286 1 272 
2 287 1 272 
2 288 1 272 
2 289 1 272 
0 290 4 1 2 282 115
0 291 4 1 2 283 119
0 292 4 1 2 284 117
0 293 4 1 2 285 121
0 294 4 1 2 286 224
0 295 4 1 2 287 231
0 296 6 1 2 277 214
0 297 3 1 2 288 228
0 298 4 1 2 278 181
0 299 6 1 2 201 279
0 300 6 1 2 280 215
0 301 4 1 2 289 226
0 302 6 1 2 281 197
0 303 4 1 2 35 294
0 304 4 1 2 295 74
0 305 6 1 2 297 112
0 306 6 1 2 300 299
0 307 4 1 2 301 86
0 308 6 1 2 303 199
0 309 6 1 2 304 219
0 310 4 1 2 305 191
0 311 6 1 2 307 188
0 312 6 1 2 309 308
0 313 4 1 2 298 310
0 314 6 1 2 302 311
0 315 6 1 2 313 296
0 316 4 1 2 314 306
0 317 4 1 2 315 312
3 318 6 0 2 316 317
2 319 1 318 
2 320 1 318 
2 321 1 318 
2 322 1 318 
2 323 1 318 
2 324 1 318 
0 325 7 1 2 85 319
0 326 7 1 2 57 320
0 327 7 1 2 79 321
0 328 5 3 1 322
0 329 7 1 2 65 323
0 330 6 1 2 52 324
0 331 4 1 2 291 325
0 332 4 1 2 292 326
0 333 4 1 2 327 293
0 334 4 1 2 329 133
0 335 6 1 2 330 44
2 336 1 328 
2 337 1 328 
2 338 1 328 
0 339 4 1 2 336 113
0 340 4 1 2 337 111
0 341 6 2 2 331 187
0 342 6 2 2 332 183
0 343 7 3 2 333 196
0 344 4 2 2 100 338
0 345 6 2 2 334 275
0 346 4 1 2 276 335
0 347 4 1 2 290 339
0 348 3 1 2 264 340
2 349 1 341 
2 350 1 341 
2 351 1 342 
2 352 1 342 
2 353 1 343 
2 354 1 343 
2 355 1 343 
2 356 1 344 
2 357 1 344 
2 358 1 345 
2 359 1 345 
0 360 3 1 2 349 353
0 361 4 1 2 274 356
0 362 6 2 2 347 220
0 363 4 2 2 348 190
0 364 5 2 1 352
0 365 4 1 2 265 357
0 366 5 2 1 359
0 367 7 2 2 365 218
2 368 1 362 
2 369 1 362 
2 370 1 363 
2 371 1 363 
2 372 1 364 
2 373 1 364 
2 374 1 366 
2 375 1 366 
0 376 4 1 2 368 370
0 377 4 1 2 372 374
0 378 5 1 1 371
0 379 4 1 2 373 355
2 380 1 367 
2 381 1 367 
0 382 4 1 2 361 376
0 383 4 1 2 354 380
0 384 6 2 2 378 350
0 385 4 1 2 381 375
0 386 6 1 2 382 360
3 387 6 0 2 385 379
2 388 1 384 
2 389 1 384 
0 390 6 1 2 386 358
0 391 6 1 2 383 388
0 392 5 1 1 389
0 393 3 1 2 387 97
3 394 6 0 2 390 351
3 395 6 0 2 377 391
0 396 6 1 2 392 369
0 397 4 1 2 393 396
3 398 4 0 2 346 397
