1 0 0 2 0
1 1 0 1 0
1 2 0 2 0
1 3 0 1 0
1 4 0 2 0
1 5 0 3 0
1 6 0 3 0
1 7 0 1 0
1 8 0 3 0
1 9 0 3 0
1 10 0 3 0
1 11 0 2 0
1 12 0 3 0
1 13 0 3 0
1 14 0 3 0
1 15 0 2 0
1 16 0 3 0
1 17 0 2 0
1 18 0 2 0
1 19 0 2 0
1 20 0 2 0
1 21 0 2 0
1 22 0 2 0
1 23 0 1 0
1 24 0 2 0
1 25 0 3 0
1 26 0 3 0
1 27 0 3 0
1 28 0 3 0
1 29 0 2 0
1 30 0 2 0
1 31 0 2 0
1 32 0 2 0
1 33 0 3 0
1 34 0 2 0
1 35 0 2 0
0 36 5 1 1 7
0 37 5 1 1 3
0 38 5 1 1 23
0 39 5 4 1 1
2 40 1 0 
2 41 1 0 
2 42 1 2 
2 43 1 2 
2 44 1 4 
2 45 1 4 
2 46 1 5 
2 47 1 5 
2 48 1 5 
2 49 1 6 
2 50 1 6 
2 51 1 6 
2 52 1 8 
2 53 1 8 
2 54 1 8 
2 55 1 9 
2 56 1 9 
2 57 1 9 
2 58 1 10 
2 59 1 10 
2 60 1 10 
2 61 1 11 
2 62 1 11 
2 63 1 12 
2 64 1 12 
2 65 1 12 
2 66 1 13 
2 67 1 13 
2 68 1 13 
2 69 1 14 
2 70 1 14 
2 71 1 14 
2 72 1 15 
2 73 1 15 
2 74 1 16 
2 75 1 16 
2 76 1 16 
2 77 1 17 
2 78 1 17 
2 79 1 18 
2 80 1 18 
2 81 1 19 
2 82 1 19 
2 83 1 20 
2 84 1 20 
2 85 1 21 
2 86 1 21 
2 87 1 22 
2 88 1 22 
2 89 1 24 
2 90 1 24 
2 91 1 25 
2 92 1 25 
2 93 1 25 
2 94 1 26 
2 95 1 26 
2 96 1 26 
2 97 1 27 
2 98 1 27 
2 99 1 27 
2 100 1 28 
2 101 1 28 
2 102 1 28 
2 103 1 29 
2 104 1 29 
2 105 1 30 
2 106 1 30 
2 107 1 31 
2 108 1 31 
2 109 1 32 
2 110 1 32 
2 111 1 33 
2 112 1 33 
2 113 1 33 
2 114 1 34 
2 115 1 34 
2 116 1 35 
2 117 1 35 
0 118 5 3 1 104
0 119 5 1 1 86
0 120 5 1 1 78
0 121 5 1 1 68
0 122 6 2 2 36 57
0 123 6 2 2 37 48
0 124 6 2 2 38 93
0 125 5 1 1 108
2 126 1 39 
2 127 1 39 
2 128 1 39 
2 129 1 39 
0 130 4 1 2 119 82
0 131 4 1 2 120 73
0 132 4 1 2 121 62
0 133 3 1 2 41 129
0 134 6 1 2 125 113
2 135 1 118 
2 136 1 118 
2 137 1 118 
2 138 1 122 
2 139 1 122 
2 140 1 123 
2 141 1 123 
2 142 1 124 
2 143 1 124 
0 144 4 1 2 99 137
0 145 7 1 3 139 141 143
0 146 4 1 4 132 131 130 144
3 147 6 0 4 134 133 145 146
2 148 1 147 
2 149 1 147 
2 150 1 147 
2 151 1 147 
2 152 1 147 
2 153 1 147 
2 154 1 147 
2 155 1 147 
2 156 1 147 
2 157 1 147 
0 158 6 1 2 97 148
0 159 6 2 2 149 142
0 160 6 2 2 61 150
0 161 6 2 2 151 138
0 162 6 2 2 152 140
0 163 6 1 2 81 153
0 164 6 1 2 72 154
0 165 7 2 2 98 155
0 166 7 3 2 40 156
0 167 6 1 2 107 157
0 168 7 2 2 158 103
0 169 6 3 2 163 85
0 170 6 3 2 164 77
0 171 6 3 2 167 112
2 172 1 159 
2 173 1 159 
2 174 1 160 
2 175 1 160 
2 176 1 161 
2 177 1 161 
2 178 1 162 
2 179 1 162 
2 180 1 165 
2 181 1 165 
2 182 1 166 
2 183 1 166 
2 184 1 166 
0 185 6 3 2 92 173
0 186 6 3 2 67 175
0 187 6 3 2 56 177
0 188 6 3 2 47 179
0 189 4 1 3 106 181 136
0 190 3 1 3 43 184 128
2 191 1 168 
2 192 1 168 
2 193 1 169 
2 194 1 169 
2 195 1 169 
2 196 1 170 
2 197 1 170 
2 198 1 170 
2 199 1 171 
2 200 1 171 
2 201 1 171 
0 202 5 1 1 193
0 203 5 1 1 196
0 204 4 1 2 116 199
0 205 3 1 3 114 117 200
0 206 4 2 2 88 195
0 207 4 2 2 80 198
0 208 3 1 2 115 201
2 209 1 185 
2 210 1 185 
2 211 1 185 
2 212 1 186 
2 213 1 186 
2 214 1 186 
2 215 1 187 
2 216 1 187 
2 217 1 187 
2 218 1 188 
2 219 1 188 
2 220 1 188 
0 221 4 1 2 53 218
0 222 4 1 2 64 215
0 223 3 1 2 75 212
0 224 3 1 2 101 209
0 225 4 1 3 95 102 210
0 226 3 1 3 50 54 219
0 227 3 1 3 59 65 216
0 228 4 1 3 70 76 213
0 229 4 1 2 96 211
0 230 4 1 2 71 214
0 231 4 1 2 60 217
0 232 4 1 2 51 220
2 233 1 206 
2 234 1 206 
2 235 1 207 
2 236 1 207 
0 237 6 1 2 224 223
0 238 6 1 2 227 226
0 239 4 1 4 232 231 230 229
0 240 4 1 3 189 234 236
0 241 4 1 4 237 222 204 221
3 242 6 0 4 208 190 240 239
2 243 1 242 
2 244 1 242 
2 245 1 242 
2 246 1 242 
2 247 1 242 
2 248 1 242 
2 249 1 242 
2 250 1 242 
2 251 1 242 
2 252 1 242 
0 253 6 1 2 94 243
0 254 6 1 2 87 244
0 255 6 1 2 58 245
0 256 6 1 2 49 246
0 257 6 1 2 79 247
0 258 6 1 2 69 248
0 259 4 1 2 241 249
0 260 5 2 1 250
0 261 6 2 2 105 251
0 262 7 2 2 42 252
0 263 4 1 4 228 238 225 259
2 264 1 260 
2 265 1 260 
2 266 1 261 
2 267 1 261 
2 268 1 262 
2 269 1 262 
0 270 4 1 2 264 235
0 271 4 1 2 265 233
0 272 5 1 1 267
0 273 3 1 4 45 269 183 127
0 274 4 1 3 270 84 197
0 275 4 1 3 271 90 194
0 276 4 1 4 272 110 180 135
0 277 4 1 3 276 275 274
3 278 6 0 4 205 273 277 263
2 279 1 278 
2 280 1 278 
2 281 1 278 
2 282 1 278 
2 283 1 278 
2 284 1 278 
2 285 1 278 
2 286 1 278 
0 287 6 1 2 109 279
0 288 6 1 2 100 280
0 289 6 1 2 89 281
0 290 6 1 2 63 282
0 291 6 1 2 52 283
0 292 6 1 2 83 284
0 293 6 1 2 74 285
0 294 7 1 2 44 286
0 295 6 2 4 288 253 91 172
0 296 6 2 3 289 254 202
0 297 6 3 4 290 255 55 176
0 298 6 3 4 291 256 46 178
0 299 6 3 3 292 257 203
0 300 6 3 4 293 258 66 174
0 301 4 1 4 294 268 182 126
2 302 1 295 
2 303 1 295 
2 304 1 296 
2 305 1 296 
2 306 1 297 
2 307 1 297 
2 308 1 297 
2 309 1 298 
2 310 1 298 
2 311 1 298 
2 312 1 299 
2 313 1 299 
2 314 1 299 
2 315 1 300 
2 316 1 300 
2 317 1 300 
0 318 5 1 1 304
0 319 6 1 4 287 302 191 266
0 320 6 2 2 303 305
3 321 6 0 4 308 311 314 317
0 322 6 1 2 318 312
2 323 1 320 
2 324 1 320 
0 325 6 1 3 319 322 315
0 326 6 1 3 323 313 316
0 327 4 1 4 321 111 324 192
0 328 6 1 2 325 306
3 329 6 0 3 326 307 310
3 330 4 0 2 301 327
3 331 6 0 2 328 309
