1 1	0 2	0
1 2	0 2	0
1 3	0 1	0
2 4	1 1
2 5	1 2
2 6	1 1
2 7	1 2
0 8	2 2	2 4 5
2 9	1 8
2 10 1 8
2 11 1 3
2 12 1 3
3 13 2 0 2 9 11
0 14 7 1 2 10 12
0 15 7 1 2 6 7
3 16 3 0 2 14 15
