1 0 0 1 0
1 1 0 2 0
1 2 0 2 0
1 3 0 1 0
1 4 0 1 0
2 5 1 1 
2 6 1 1 
2 7 1 2 
2 8 1 2 
0 9 4 1 2 4 5
0 10 6 2 2 3 7
0 11 6 1 2 0 8
2 12 1 10 
2 13 1 10 
0 14 5 1 1 12
0 15 6 1 2 6 13
3 16 4 0 2 14 9
3 17 6 0 2 11 15
