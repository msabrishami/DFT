1 N1 0 5 0
1 N8 0 2 0
1 N13 0 3 0
1 N17 0 5 0
1 N26 0 1 0
1 N29 0 3 0
1 N36 0 4 0
1 N42 0 4 0
1 N51 0 2 0
1 N55 0 3 0
1 N59 0 4 0
1 N68 0 1 0
1 N72 0 1 0
1 N73 0 1 0
1 N74 0 1 0
1 N75 0 2 0
1 N80 0 2 0
1 N85 0 1 0
1 N86 0 1 0
1 N87 0 1 0
1 N88 0 1 0
1 N89 0 1 0
1 N90 0 1 0
1 N91 0 3 0
1 N96 0 3 0
1 N101 0 1 0
1 N106 0 2 0
1 N111 0 2 0
1 N116 0 4 0
1 N121 0 4 0
1 N126 0 3 0
1 N130 0 5 0
1 N135 0 3 0
1 N138 0 2 0
1 N143 0 2 0
1 N146 0 2 0
1 N149 0 2 0
1 N152 0 1 0
1 N153 0 2 0
1 N156 0 1 0
1 N159 0 3 0
1 N165 0 4 0
1 N171 0 5 0
1 N177 0 4 0
1 N183 0 4 0
1 N189 0 4 0
1 N195 0 5 0
1 N201 0 5 0
1 N207 0 3 0
1 N210 0 4 0
1 N219 0 8 0
1 N228 0 3 0
1 N237 0 8 0
1 N246 0 6 0
1 N255 0 3 0
1 N259 0 1 0
1 N260 0 1 0
1 N261 0 3 0
1 N267 0 1 0
1 N268 0 2 0
0 n601 7 1 2 N73 N72
0 n450 5 4 1 N101
0 n721 3 2 2 N87 N88
3 N391 7 0 2 N86 N85
0 n740 5 1 1 N26
2 N1-1 1 N1 
2 N1-2 1 N1 
2 N1-3 1 N1 
2 N1-4 1 N1 
2 N1-5 1 N1 
2 N8-1 1 N8 
2 N8-2 1 N8 
2 N13-1 1 N13 
2 N13-2 1 N13 
2 N13-3 1 N13 
2 N17-1 1 N17 
2 N17-2 1 N17 
2 N17-3 1 N17 
2 N17-4 1 N17 
2 N17-5 1 N17 
2 N29-1 1 N29 
2 N29-2 1 N29 
2 N29-3 1 N29 
2 N36-1 1 N36 
2 N36-2 1 N36 
2 N36-3 1 N36 
2 N36-4 1 N36 
2 N42-1 1 N42 
2 N42-2 1 N42 
2 N42-3 1 N42 
2 N42-4 1 N42 
2 N51-1 1 N51 
2 N51-2 1 N51 
2 N55-1 1 N55 
2 N55-2 1 N55 
2 N55-3 1 N55 
2 N59-1 1 N59 
2 N59-2 1 N59 
2 N59-3 1 N59 
2 N59-4 1 N59 
2 N75-1 1 N75 
2 N75-2 1 N75 
2 N80-1 1 N80 
2 N80-2 1 N80 
2 N91-1 1 N91 
2 N91-2 1 N91 
2 N91-3 1 N91 
2 N96-1 1 N96 
2 N96-2 1 N96 
2 N96-3 1 N96 
2 N106-1 1 N106 
2 N106-2 1 N106 
2 N111-1 1 N111 
2 N111-2 1 N111 
2 N116-1 1 N116 
2 N116-2 1 N116 
2 N116-3 1 N116 
2 N116-4 1 N116 
2 N121-1 1 N121 
2 N121-2 1 N121 
2 N121-3 1 N121 
2 N121-4 1 N121 
2 N126-1 1 N126 
2 N126-2 1 N126 
2 N126-3 1 N126 
2 N130-1 1 N130 
2 N130-2 1 N130 
2 N130-3 1 N130 
2 N130-4 1 N130 
2 N130-5 1 N130 
2 N135-1 1 N135 
2 N135-2 1 N135 
2 N135-3 1 N135 
2 N138-1 1 N138 
2 N138-2 1 N138 
2 N143-1 1 N143 
2 N143-2 1 N143 
2 N146-1 1 N146 
2 N146-2 1 N146 
2 N149-1 1 N149 
2 N149-2 1 N149 
2 N153-1 1 N153 
2 N153-2 1 N153 
2 N159-1 1 N159 
2 N159-2 1 N159 
2 N159-3 1 N159 
2 N165-1 1 N165 
2 N165-2 1 N165 
2 N165-3 1 N165 
2 N165-4 1 N165 
2 N171-1 1 N171 
2 N171-2 1 N171 
2 N171-3 1 N171 
2 N171-4 1 N171 
2 N171-5 1 N171 
2 N177-1 1 N177 
2 N177-2 1 N177 
2 N177-3 1 N177 
2 N177-4 1 N177 
2 N183-1 1 N183 
2 N183-2 1 N183 
2 N183-3 1 N183 
2 N183-4 1 N183 
2 N189-1 1 N189 
2 N189-2 1 N189 
2 N189-3 1 N189 
2 N189-4 1 N189 
2 N195-1 1 N195 
2 N195-2 1 N195 
2 N195-3 1 N195 
2 N195-4 1 N195 
2 N195-5 1 N195 
2 N201-1 1 N201 
2 N201-2 1 N201 
2 N201-3 1 N201 
2 N201-4 1 N201 
2 N201-5 1 N201 
2 N207-1 1 N207 
2 N207-2 1 N207 
2 N207-3 1 N207 
2 N210-1 1 N210 
2 N210-2 1 N210 
2 N210-3 1 N210 
2 N210-4 1 N210 
2 N219-1 1 N219 
2 N219-2 1 N219 
2 N219-3 1 N219 
2 N219-4 1 N219 
2 N219-5 1 N219 
2 N219-6 1 N219 
2 N219-7 1 N219 
2 N219-8 1 N219 
2 N228-1 1 N228 
2 N228-2 1 N228 
2 N228-3 1 N228 
2 N237-1 1 N237 
2 N237-2 1 N237 
2 N237-3 1 N237 
2 N237-4 1 N237 
2 N237-5 1 N237 
2 N237-6 1 N237 
2 N237-7 1 N237 
2 N237-8 1 N237 
2 N246-1 1 N246 
2 N246-2 1 N246 
2 N246-3 1 N246 
2 N246-4 1 N246 
2 N246-5 1 N246 
2 N246-6 1 N246 
2 N255-1 1 N255 
2 N255-2 1 N255 
2 N255-3 1 N255 
2 N261-1 1 N261 
2 N261-2 1 N261 
2 N261-3 1 N261 
2 N268-1 1 N268 
2 N268-2 1 N268 
0 n426 7 1 2 N210-1 N268-1
0 n444 5 1 1 N149-1
0 n454 5 1 1 N146-1
0 n463 5 1 1 N143-1
0 n448 5 3 1 N138-1
0 n492 5 1 1 N153-1
0 n499 7 1 2 N152 N138-2
0 n515 6 1 2 N116-1 N210-2
0 n514 6 1 2 N260 N255-1
0 n530 6 1 2 N259 N255-2
0 n523 5 2 1 N219-6
0 n387 5 5 1 N210-3
0 n596 5 1 1 N261-2
0 n604 6 1 2 N42-1 N59-1
0 n410 5 3 1 N246-6
0 n609 6 1 2 N121-1 N210-4
0 n608 6 1 2 N267 N255-3
0 n386 5 6 1 N228-3
0 n494 7 3 2 N156 N59-2
0 n457 5 2 1 N51-1
0 n447 5 3 1 N17-3
0 n459 5 3 1 N159-2
0 n434 5 2 1 N165-4
0 n378 5 3 1 N171-4
0 n483 5 4 1 N177-4
0 n578 5 4 1 N183-3
0 n547 5 4 1 N189-4
0 n511 5 3 1 N195-5
0 n614 5 3 1 N201-4
0 n648 5 2 1 N207-3
0 n571 5 3 1 N121-4
0 n500 5 3 1 N106-1
0 n533 5 3 1 N111-2
0 n575 5 3 1 N116-3
0 n712 5 2 1 N130-5
0 n408 5 4 1 N91-2
0 n388 5 4 1 N96-3
0 n619 5 3 1 N126-2
0 n688 5 2 1 N135-3
0 n725 6 1 2 N1-3 N55-3
0 n466 5 3 1 N8-1
0 n723 7 1 2 N68 N13-1
0 n633 5 4 1 N59-3
0 n729 5 2 1 N80-1
0 n632 5 2 1 N75-1
0 n731 7 1 2 N13-2 N17-4
0 n734 6 1 2 N8-2 N13-3
0 n733 6 1 2 N1-4 N17-5
0 n637 5 3 1 N29-1
0 n737 6 1 2 N29-2 N80-2
0 n736 5 1 1 N36-4
0 n738 6 1 2 N29-3 N75-2
0 n626 5 4 1 N42-4
0 n739 5 1 1 N1-5
2 n450-1 1 n450 
2 n450-2 1 n450 
2 n450-3 1 n450 
2 n450-4 1 n450 
2 n721-1 1 n721 
2 n721-2 1 n721 
0 n513 6 1 2 n514 n515
0 n607 6 1 2 n608 n609
3 N450 7 0 2 N89 n721-1
3 N423 7 0 2 N90 n721-2
3 N418 4 0 2 n733 n734
3 N389 4 0 2 n736 n737
0 n732 4 2 2 n739 n740
2 n448-1 1 n448 
2 n448-2 1 n448 
2 n448-3 1 n448 
2 n523-1 1 n523 
2 n523-2 1 n523 
2 n387-1 1 n387 
2 n387-2 1 n387 
2 n387-3 1 n387 
2 n387-4 1 n387 
2 n387-5 1 n387 
2 n410-1 1 n410 
2 n410-2 1 n410 
2 n410-3 1 n410 
2 n386-1 1 n386 
2 n386-2 1 n386 
2 n386-3 1 n386 
2 n386-4 1 n386 
2 n386-5 1 n386 
2 n386-6 1 n386 
2 n494-1 1 n494 
2 n494-2 1 n494 
2 n494-3 1 n494 
2 n457-1 1 n457 
2 n457-2 1 n457 
2 n447-1 1 n447 
2 n447-2 1 n447 
2 n447-3 1 n447 
2 n459-1 1 n459 
2 n459-2 1 n459 
2 n459-3 1 n459 
2 n434-1 1 n434 
2 n434-2 1 n434 
2 n378-1 1 n378 
2 n378-2 1 n378 
2 n378-3 1 n378 
2 n483-1 1 n483 
2 n483-2 1 n483 
2 n483-3 1 n483 
2 n483-4 1 n483 
2 n578-1 1 n578 
2 n578-2 1 n578 
2 n578-3 1 n578 
2 n578-4 1 n578 
2 n547-1 1 n547 
2 n547-2 1 n547 
2 n547-3 1 n547 
2 n547-4 1 n547 
2 n511-1 1 n511 
2 n511-2 1 n511 
2 n511-3 1 n511 
2 n614-1 1 n614 
2 n614-2 1 n614 
2 n614-3 1 n614 
2 n648-1 1 n648 
2 n648-2 1 n648 
2 n571-1 1 n571 
2 n571-2 1 n571 
2 n571-3 1 n571 
2 n500-1 1 n500 
2 n500-2 1 n500 
2 n500-3 1 n500 
2 n533-1 1 n533 
2 n533-2 1 n533 
2 n533-3 1 n533 
2 n575-1 1 n575 
2 n575-2 1 n575 
2 n575-3 1 n575 
2 n712-1 1 n712 
2 n712-2 1 n712 
2 n408-1 1 n408 
2 n408-2 1 n408 
2 n408-3 1 n408 
2 n408-4 1 n408 
2 n388-1 1 n388 
2 n388-2 1 n388 
2 n388-3 1 n388 
2 n388-4 1 n388 
2 n619-1 1 n619 
2 n619-2 1 n619 
2 n619-3 1 n619 
2 n688-1 1 n688 
2 n688-2 1 n688 
2 n466-1 1 n466 
2 n466-2 1 n466 
2 n466-3 1 n466 
2 n633-1 1 n633 
2 n633-2 1 n633 
2 n633-3 1 n633 
2 n633-4 1 n633 
2 n729-1 1 n729 
2 n729-2 1 n729 
2 n632-1 1 n632 
2 n632-2 1 n632 
2 n637-1 1 n637 
2 n637-2 1 n637 
2 n637-3 1 n637 
2 n626-1 1 n626 
2 n626-2 1 n626 
2 n626-3 1 n626 
2 n626-4 1 n626 
0 n380 4 1 2 n387-1 n388-1
0 n407 4 1 2 n387-2 n408-1
0 n446 4 1 2 n448-1 n447-1
0 n456 4 1 2 n448-2 n457-1
0 n465 4 1 2 n448-3 n466-1
0 n485 4 1 2 n387-3 n450-2
0 n532 4 1 2 n387-4 n533-1
0 n580 4 1 2 n387-5 n500-2
0 n625 4 1 2 N42-2 n447-2
0 n624 4 1 2 N17-2 n626-1
0 n631 4 1 2 n633-1 n632-1
0 n627 4 1 2 n447-3 n466-2
0 n636 4 1 2 N268-2 n637-1
0 n647 6 1 2 N207-1 n614-2
0 n646 6 1 2 N201-3 n648-1
0 n658 6 1 2 N165-3 n459-3
0 n657 6 1 2 N159-3 n434-2
0 n667 6 1 2 N189-2 n578-3
0 n666 6 1 2 N183-2 n547-3
0 n669 4 1 2 N177-2 n378-2
0 n668 4 1 2 N171-3 n483-3
0 n673 6 1 2 N177-3 n378-3
0 n672 6 1 2 N171-5 n483-4
0 n675 4 1 2 N189-3 n578-4
0 n674 4 1 2 N183-4 n547-4
0 n677 4 1 2 N207-2 n614-3
0 n676 4 1 2 N201-5 n648-2
0 n687 6 1 2 N135-1 n619-2
0 n686 6 1 2 N126-1 n688-1
0 n705 6 1 2 N111-1 n500-3
0 n704 6 1 2 N106-2 n533-3
0 n709 6 1 2 N96-1 n408-3
0 n708 6 1 2 N91-1 n388-3
0 n711 4 1 2 N130-3 n575-2
0 n710 4 1 2 N116-2 n712-1
0 n716 6 1 2 N130-4 n575-3
0 n715 6 1 2 N116-4 n712-2
0 n718 4 1 2 N96-2 n408-4
0 n717 4 1 2 N91-3 n388-4
0 n720 4 1 2 N135-2 n619-3
0 n719 4 1 2 N126-3 n688-2
0 n724 4 1 2 n725 n466-3
0 n727 4 1 2 n633-3 n626-2
0 n728 4 1 2 n633-4 n729-1
0 n635 4 2 2 n729-2 n632-2
0 n735 4 1 2 n637-3 n626-3
3 N388 4 0 2 n738 n626-4
2 n732-1 1 n732 
2 n732-2 1 n732 
0 n623 4 1 2 n624 n625
0 n630 6 1 2 n631 N42-3
0 n640 6 1 2 n646 n647
0 n655 6 2 2 n657 n658
0 n665 6 1 2 n666 n667
0 n664 4 1 2 n668 n669
0 n671 6 1 2 n672 n673
0 n670 4 1 2 n674 n675
0 n649 4 1 2 n676 n677
0 n680 6 1 2 n686 n687
0 n703 6 2 2 n704 n705
0 n707 6 1 2 n708 n709
0 n706 4 1 2 n710 n711
0 n714 6 1 2 n715 n716
0 n713 4 1 2 n717 n718
0 n689 4 1 2 n719 n720
0 n603 6 3 2 n723 n724
3 N422 6 0 2 n727 N36-1
3 N421 6 0 2 n728 N36-2
0 n726 7 2 2 n731 n732-1
0 n730 6 2 2 n735 N36-3
0 n495 6 4 2 N51-2 n732-2
2 n635-1 1 n635 
2 n635-2 1 n635 
0 n629 6 1 2 n630 N1-2
0 n497 6 2 2 n636 n635-1
0 n663 6 1 2 n664 n665
0 n662 6 1 2 n670 n671
0 n697 6 2 2 n706 n707
0 n698 6 2 2 n713 n714
3 N420 6 0 2 N59-4 n635-2
2 n655-1 1 n655 
2 n655-2 1 n655 
2 n703-1 1 n703 
2 n703-2 1 n703 
2 n603-1 1 n603 
2 n603-2 1 n603 
2 n603-3 1 n603 
2 n726-1 1 n726 
2 n726-2 1 n726 
2 n730-1 1 n730 
2 n730-2 1 n730 
2 n495-1 1 n495 
2 n495-2 1 n495 
2 n495-3 1 n495 
2 n495-4 1 n495 
0 n493 4 1 2 n494-1 n495-1
0 n602 4 1 2 n604 n603-1
0 n622 4 1 2 n623 n495-2
0 n628 4 1 2 n629 n457-2
0 n661 6 2 2 n662 n663
0 n699 4 2 2 n450-3 n703-1
0 n700 7 2 2 n450-4 n703-2
0 n722 4 1 2 n603-2 n633-2
3 N448 4 0 2 n603-3 n637-2
3 N419 6 0 2 n726-2 n730-1
3 N390 5 0 1 n730-2
3 N447 5 0 1 n495-4
2 n497-1 1 n497 
2 n497-2 1 n497 
2 n697-1 1 n697 
2 n697-2 1 n697 
2 n698-1 1 n698 
2 n698-2 1 n698 
0 n443 6 4 2 n493 N55-1
0 n379 6 4 2 n601 n602
0 n496 6 2 2 N447 N17-1
0 n621 6 1 2 n622 n494-3
0 n620 6 1 2 n627 n628
0 n634 4 1 2 n497-2 n495-3
0 n696 6 1 2 n697-1 n698-1
0 n701 7 1 2 n697-2 n698-2
3 N449 7 0 2 n722 N74
3 N446 6 0 2 N390 n726-1
2 n661-1 1 n661 
2 n661-2 1 n661 
2 n699-1 1 n699 
2 n699-2 1 n699 
2 n700-1 1 n700 
2 n700-2 1 n700 
0 n449 7 8 2 n620 n621
0 n569 7 4 2 n634 N55-2
0 n660 6 1 2 N130-1 n661-1
0 n659 3 1 2 N130-2 n661-2
0 n695 4 1 2 n699-1 n700-1
0 n702 3 1 2 n699-2 n700-2
2 n443-1 1 n443 
2 n443-2 1 n443 
2 n443-3 1 n443 
2 n443-4 1 n443 
2 n379-1 1 n379 
2 n379-2 1 n379 
2 n379-3 1 n379 
2 n379-4 1 n379 
2 n496-1 1 n496 
2 n496-2 1 n496 
0 n361 4 1 2 n379-1 n378-1
0 n442 4 1 2 n444 n443-1
0 n453 4 1 2 n454 n443-2
0 n462 4 1 2 n463 n443-3
0 n491 4 1 2 n492 n443-4
0 n441 4 4 2 n496-1 n497-1
0 n503 4 1 2 n379-3 n511-1
0 n431 5 5 1 n379-4
0 n617 3 1 2 n496-2 n494-2
0 n656 7 2 2 n659 n660
0 n694 6 1 2 n695 n696
0 n693 6 1 2 n701 n702
2 n449-1 1 n449 
2 n449-2 1 n449 
2 n449-3 1 n449 
2 n449-4 1 n449 
2 n449-5 1 n449 
2 n449-6 1 n449 
2 n449-7 1 n449 
2 n449-8 1 n449 
2 n569-1 1 n569 
2 n569-2 1 n569 
2 n569-3 1 n569 
2 n569-4 1 n569 
0 n445 4 1 2 n449-1 n450-1
0 n455 4 1 2 n449-2 n388-2
0 n464 4 1 2 n449-3 n408-2
0 n498 4 1 2 n449-4 n500-1
0 n570 4 1 2 n449-5 n571-1
0 n574 4 1 2 n449-6 n575-1
0 n586 4 1 2 n449-7 n533-2
0 n568 6 4 2 n617 N1-1
0 n618 4 1 2 n449-8 n619-1
0 n684 6 3 2 n693 n694
2 n441-1 1 n441 
2 n441-2 1 n441 
2 n441-3 1 n441 
2 n441-4 1 n441 
2 n431-1 1 n431 
2 n431-2 1 n431 
2 n431-3 1 n431 
2 n431-4 1 n431 
2 n431-5 1 n431 
2 n656-1 1 n656 
2 n656-2 1 n656 
0 n428 6 1 2 N159-1 n431-1
0 n440 4 1 2 n442 n441-1
0 n439 4 1 2 n445 n446
0 n452 4 1 2 n453 n441-2
0 n451 4 1 2 n455 n456
0 n461 4 1 2 n462 n441-3
0 n460 4 1 2 n464 n465
0 n490 4 1 2 n491 n441-4
0 n489 4 1 2 n498 n499
0 n487 6 1 2 N177-1 n431-2
0 n566 4 1 2 n570 n569-1
0 n572 4 1 2 n574 n569-2
0 n584 4 1 2 n586 n569-3
0 n582 6 1 2 N183-1 n431-4
0 n591 6 1 2 N201-1 n431-5
0 n615 4 1 2 n618 n569-4
0 n654 6 1 2 n655-1 n656-1
0 n653 3 1 2 n655-2 n656-2
2 n568-1 1 n568 
2 n568-2 1 n568 
2 n568-3 1 n568 
2 n568-4 1 n568 
2 n684-1 1 n684 
2 n684-2 1 n684 
2 n684-3 1 n684 
0 n377 6 3 2 n439 n440
0 n403 6 3 2 n451 n452
0 n430 6 2 2 n460 n461
0 n484 6 2 2 n489 n490
0 n567 6 1 2 N149-2 n568-1
0 n573 6 1 2 N146-2 n568-2
0 n585 6 1 2 N143-2 n568-3
0 n616 6 1 2 N153-2 n568-4
0 n645 6 3 2 n653 n654
0 n683 6 1 2 N121-2 n684-1
0 n692 4 1 2 N121-3 n684-2
0 n685 5 2 1 n684-3
0 n510 6 3 2 n566 n567
0 n549 6 3 2 n572 n573
0 n579 6 2 2 n584 n585
0 n613 6 2 2 n615 n616
2 n377-1 1 n377 
2 n377-2 1 n377 
2 n377-3 1 n377 
2 n403-1 1 n403 
2 n403-2 1 n403 
2 n403-3 1 n403 
2 n430-1 1 n430 
2 n430-2 1 n430 
2 n484-1 1 n484 
2 n484-2 1 n484 
2 n645-1 1 n645 
2 n645-2 1 n645 
2 n645-3 1 n645 
2 n685-1 1 n685 
2 n685-2 1 n685 
0 n363 6 1 2 N246-1 n377-1
0 n402 6 1 2 N237-2 n403-1
0 n429 6 1 2 N246-2 n430-1
0 n409 5 2 1 n403-2
0 n385 6 3 2 N171-1 n377-2
0 n374 4 4 2 N171-2 n377-3
0 n404 6 2 2 N165-2 n403-3
0 n458 5 2 1 n430-2
0 n482 5 2 1 n484-1
0 n488 6 1 2 N246-3 n484-2
0 n642 6 1 2 n645-1 n511-2
0 n644 5 2 1 n645-2
0 n651 4 1 2 n645-3 n511-3
0 n682 6 1 2 n571-2 n685-1
0 n691 4 1 2 n571-3 n685-2
2 n510-1 1 n510 
2 n510-2 1 n510 
2 n510-3 1 n510 
2 n549-1 1 n549 
2 n549-2 1 n549 
2 n549-3 1 n549 
2 n579-1 1 n579 
2 n579-2 1 n579 
2 n613-1 1 n613 
2 n613-2 1 n613 
0 n401 6 1 2 n402 n379-2
0 n427 6 1 2 n428 n429
0 n486 6 1 2 n487 n488
0 n505 6 1 2 N246-4 n510-1
0 n548 7 1 2 N237-6 n549-1
0 n534 5 2 1 n549-2
0 n520 4 3 2 N195-1 n510-2
0 n519 6 3 2 N195-2 n510-3
0 n544 6 2 2 N189-1 n549-3
0 n577 5 2 1 n579-1
0 n583 6 1 2 N246-5 n579-2
0 n598 4 3 2 N201-2 n613-1
0 n605 5 2 1 n613-2
0 n681 6 1 2 n682 n683
0 n690 4 1 2 n691 n692
2 n409-1 1 n409 
2 n409-2 1 n409 
2 n385-1 1 n385 
2 n385-2 1 n385 
2 n385-3 1 n385 
2 n374-1 1 n374 
2 n374-2 1 n374 
2 n374-3 1 n374 
2 n374-4 1 n374 
2 n404-1 1 n404 
2 n404-2 1 n404 
2 n458-1 1 n458 
2 n458-2 1 n458 
2 n482-1 1 n482 
2 n482-2 1 n482 
2 n644-1 1 n644 
2 n644-2 1 n644 
0 n384 4 1 2 n374-2 n386-1
0 n375 5 3 1 n385-2
0 n393 6 1 2 n401 N165-1
0 n406 4 1 2 n409-1 n410-1
0 n411 4 1 2 n426 n427
0 n405 6 2 2 n409-2 n434-1
0 n425 6 2 2 n458-1 n459-1
0 n423 4 2 2 n458-2 n459-2
0 n372 6 3 2 n482-1 n483-1
0 n481 4 2 2 n482-2 n483-2
0 n467 4 1 2 n485 n486
0 n546 4 1 2 n548 n431-3
0 n581 6 1 2 n582 n583
0 n643 6 1 2 N195-3 n644-1
0 n652 4 1 2 N195-4 n644-2
0 n679 6 1 2 n680 n681
0 n678 6 1 2 n689 n690
2 n534-1 1 n534 
2 n534-2 1 n534 
2 n520-1 1 n520 
2 n520-2 1 n520 
2 n520-3 1 n520 
2 n519-1 1 n519 
2 n519-2 1 n519 
2 n519-3 1 n519 
2 n544-1 1 n544 
2 n544-2 1 n544 
2 n577-1 1 n577 
2 n577-2 1 n577 
2 n598-1 1 n598 
2 n598-2 1 n598 
2 n598-3 1 n598 
2 n605-1 1 n605 
2 n605-2 1 n605 
0 n383 6 1 2 n384 n385-1
0 n389 4 1 2 n406 n407
0 n526 5 2 1 n519-2
0 n531 4 1 2 n534-1 n410-2
0 n538 4 1 2 n546 n547-1
0 n545 6 2 2 n534-2 n547-2
0 n479 6 2 2 n577-1 n578-1
0 n576 4 2 2 n577-2 n578-2
0 n550 4 1 2 n580 n581
0 n565 5 2 1 n598-1
0 n589 4 1 2 n410-3 n605-1
0 n612 4 1 2 n386-6 n598-3
0 n600 4 3 2 n605-2 n614-1
0 n641 6 1 2 n642 n643
0 n650 4 1 2 n651 n652
3 N767 6 0 2 n678 n679
2 n375-1 1 n375 
2 n375-2 1 n375 
2 n375-3 1 n375 
2 n405-1 1 n405 
2 n405-2 1 n405 
2 n425-1 1 n425 
2 n425-2 1 n425 
2 n423-1 1 n423 
2 n423-2 1 n423 
2 n372-1 1 n372 
2 n372-2 1 n372 
2 n372-3 1 n372 
2 n481-1 1 n481 
2 n481-2 1 n481 
0 n368 4 1 2 n375-1 n374-1
0 n382 6 1 2 N237-1 n375-3
0 n400 6 2 2 n405-1 n404-1
0 n415 6 1 2 N237-3 n423-1
0 n424 5 2 1 n423-2
0 n471 6 1 2 N237-4 n481-1
0 n371 5 3 1 n481-2
0 n529 4 1 2 n531 n532
0 n639 6 1 2 n640 n641
0 n638 6 1 2 n649 n650
2 n526-1 1 n526 
2 n526-2 1 n526 
2 n545-1 1 n545 
2 n545-2 1 n545 
2 n479-1 1 n479 
2 n479-2 1 n479 
2 n576-1 1 n576 
2 n576-2 1 n576 
2 n565-1 1 n565 
2 n565-2 1 n565 
2 n600-1 1 n600 
2 n600-2 1 n600 
2 n600-3 1 n600 
0 n381 6 1 2 n382 n383
0 n524 4 1 2 n526-1 n520-2
0 n516 6 1 2 N237-5 n526-2
0 n528 6 1 2 n529 n530
0 n537 7 3 2 n545-1 n544-1
0 n564 6 1 2 N261-1 n565-1
0 n554 6 1 2 N237-7 n576-1
0 n477 5 2 1 n576-2
0 n599 4 1 2 n598-2 n600-1
0 n563 5 3 1 n600-2
0 n610 6 1 2 N237-8 n600-3
3 N768 6 0 2 n638 n639
2 n400-1 1 n400 
2 n400-2 1 n400 
2 n424-1 1 n424 
2 n424-2 1 n424 
2 n371-1 1 n371 
2 n371-2 1 n371 
2 n371-3 1 n371 
0 n359 4 1 2 n380 n381
0 n398 5 2 1 n400-1
0 n391 4 1 2 n400-2 n386-2
0 n422 6 2 2 n425-1 n424-1
0 n436 3 1 2 n374-3 n371-2
0 n476 6 3 2 n372-3 n371-3
0 n594 4 1 2 n599 N261-3
2 n537-1 1 n537 
2 n537-2 1 n537 
2 n537-3 1 n537 
2 n477-1 1 n477 
2 n477-2 1 n477 
2 n563-1 1 n563 
2 n563-2 1 n563 
2 n563-3 1 n563 
0 n536 6 1 2 N228-2 n537-1
0 n525 6 2 2 n564 n563-1
0 n560 6 3 2 n479-2 n477-2
0 n597 6 1 2 n565-2 n563-2
0 n611 6 1 2 n612 n563-3
2 n398-1 1 n398 
2 n398-2 1 n398 
2 n422-1 1 n422 
2 n422-2 1 n422 
2 n476-1 1 n476 
2 n476-2 1 n476 
2 n476-3 1 n476 
0 n420 5 2 1 n422-1
0 n413 4 1 2 n422-2 n386-3
0 n469 4 1 2 n476-3 n386-4
0 n595 4 1 2 n596 n597
0 n606 6 1 2 n610 n611
2 n525-1 1 n525 
2 n525-2 1 n525 
2 n560-1 1 n560 
2 n560-2 1 n560 
2 n560-3 1 n560 
0 n508 7 2 2 n524 n525-1
0 n509 5 2 1 n525-2
0 n552 4 1 2 n560-3 n386-5
0 n593 4 1 2 n594 n595
0 n587 4 1 2 n606 n607
2 n420-1 1 n420 
2 n420-2 1 n420 
0 n592 6 1 2 n593 N219-8
2 n508-1 1 n508 
2 n508-2 1 n508 
2 n509-1 1 n509 
2 n509-2 1 n509 
0 n507 4 1 2 n508-1 n509-1
0 n522 4 1 2 n508-2 n523-1
0 n562 3 1 2 n520-3 n509-2
0 n590 6 1 2 n591 n592
0 n506 6 1 2 n507 N219-5
0 n521 4 1 2 n522 N228-1
0 n543 6 3 2 n562 n519-3
0 n588 4 1 2 n589 n590
0 n504 6 1 2 n505 n506
0 n518 4 1 2 n521 n520-1
3 N850 6 0 2 n587 n588
2 n543-1 1 n543 
2 n543-2 1 n543 
2 n543-3 1 n543 
0 n502 4 1 2 n503 n504
0 n517 6 1 2 n518 n519-1
0 n542 6 1 2 n537-2 n543-1
0 n541 3 1 2 n537-3 n543-2
0 n561 6 1 2 n545-2 n543-3
0 n512 6 1 2 n516 n517
0 n540 6 1 2 n541 n542
0 n480 6 2 2 n561 n544-2
0 n501 4 1 2 n512 n513
0 n539 4 1 2 n540 n523-2
2 n480-1 1 n480 
2 n480-2 1 n480 
0 n478 6 1 2 n480-1 n479-1
3 N865 6 0 2 n501 n502
0 n535 4 1 2 n538 n539
0 n559 5 2 1 n480-2
0 n373 6 2 2 n478 n477-1
0 n527 6 1 2 n535 n536
2 n559-1 1 n559 
2 n559-2 1 n559 
3 N864 3 0 2 n527 n528
0 n558 4 1 2 n559-1 n560-1
0 n557 7 1 2 n559-2 n560-2
2 n373-1 1 n373 
2 n373-2 1 n373 
0 n370 6 1 2 n373-1 n372-1
0 n438 5 3 1 n373-2
0 n556 4 1 2 n557 n558
0 n369 6 1 2 n370 n371-1
0 n555 6 1 2 n556 N219-7
2 n438-1 1 n438 
2 n438-2 1 n438 
2 n438-3 1 n438 
0 n367 4 1 2 n368 n369
0 n437 4 1 2 n374-4 n438-1
0 n475 4 1 2 n438-2 n476-1
0 n474 7 1 2 n438-3 n476-2
0 n553 6 1 2 n554 n555
0 n435 6 1 2 n437 n372-2
0 n473 4 1 2 n474 n475
0 n551 4 1 2 n552 n553
0 n376 7 2 2 n435 n436
0 n472 6 1 2 n473 N219-4
3 N863 6 0 2 n550 n551
0 n470 6 1 2 n471 n472
2 n376-1 1 n376 
2 n376-2 1 n376 
0 n366 4 1 2 n375-2 n376-1
0 n399 6 3 2 n385-3 n376-2
0 n468 4 1 2 n469 n470
0 n365 4 1 2 n366 n367
3 N874 6 0 2 n467 n468
2 n399-1 1 n399 
2 n399-2 1 n399 
2 n399-3 1 n399 
0 n364 6 1 2 n365 N219-1
0 n397 4 1 2 n398-1 n399-1
0 n396 7 1 2 n398-2 n399-2
0 n433 6 1 2 n405-2 n399-3
0 n362 6 1 2 n363 n364
0 n395 4 1 2 n396 n397
0 n421 6 3 2 n433 n404-2
0 n360 4 1 2 n361 n362
0 n394 6 1 2 n395 N219-2
2 n421-1 1 n421 
2 n421-2 1 n421 
2 n421-3 1 n421 
3 N880 6 0 2 n359 n360
0 n392 6 1 2 n393 n394
0 n419 4 1 2 n420-1 n421-1
0 n418 7 1 2 n420-2 n421-2
0 n432 6 1 2 n421-3 n425-2
0 n390 4 1 2 n391 n392
0 n417 4 1 2 n418 n419
3 N866 6 0 2 n432 n424-2
3 N879 6 0 2 n389 n390
0 n416 6 1 2 n417 N219-3
0 n414 6 1 2 n415 n416
0 n412 4 1 2 n413 n414
3 N878 6 0 2 n411 n412
