1 1 0 11 0 
2 2 1 1  
2 3 1 1  
2 4 1 1  
2 5 1 1  
2 6 1 1  
2 7 1 1  
2 8 1 1  
2 9 1 1  
2 10 1 1  
2 11 1 1  
2 12 1 1  
1 13 0 6 0 
2 14 1 13  
2 15 1 13  
2 16 1 13  
2 17 1 13  
2 18 1 13  
2 19 1 13  
1 20 0 12 0 
2 21 1 20  
2 22 1 20  
2 23 1 20  
2 24 1 20  
2 25 1 20  
2 26 1 20  
2 27 1 20  
2 28 1 20  
2 29 1 20  
2 30 1 20  
2 31 1 20  
2 32 1 20  
1 33 0 7 0 
2 34 1 33  
2 35 1 33  
2 36 1 33  
2 37 1 33  
2 38 1 33  
2 39 1 33  
2 40 1 33  
1 41 0 3 0 
2 42 1 41  
2 43 1 41  
2 44 1 41  
1 45 0 4 0 
2 46 1 45  
2 47 1 45  
2 48 1 45  
2 49 1 45  
1 50 0 7 0 
2 51 1 50  
2 52 1 50  
2 53 1 50  
2 54 1 50  
2 55 1 50  
2 56 1 50  
2 57 1 50  
1 58 0 9 0 
2 59 1 58  
2 60 1 58  
2 61 1 58  
2 62 1 58  
2 63 1 58  
2 64 1 58  
2 65 1 58  
2 66 1 58  
2 67 1 58  
1 68 0 8 0 
2 69 1 68  
2 70 1 68  
2 71 1 68  
2 72 1 68  
2 73 1 68  
2 74 1 68  
2 75 1 68  
2 76 1 68  
1 77 0 9 0 
2 78 1 77  
2 79 1 77  
2 80 1 77  
2 81 1 77  
2 82 1 77  
2 83 1 77  
2 84 1 77  
2 85 1 77  
2 86 1 77  
1 87 0 9 0 
2 88 1 87  
2 89 1 87  
2 90 1 87  
2 91 1 87  
2 92 1 87  
2 93 1 87  
2 94 1 87  
2 95 1 87  
2 96 1 87  
1 97 0 9 0 
2 98 1 97  
2 99 1 97  
2 100 1 97  
2 101 1 97  
2 102 1 97  
2 103 1 97  
2 104 1 97  
2 105 1 97  
2 106 1 97  
1 107 0 8 0 
2 108 1 107  
2 109 1 107  
2 110 1 107  
2 111 1 107  
2 112 1 107  
2 113 1 107  
2 114 1 107  
2 115 1 107  
1 116 0 7 0 
2 117 1 116  
2 118 1 116  
2 119 1 116  
2 120 1 116  
2 121 1 116  
2 122 1 116  
2 123 1 116  
1 124 0 1 0 
1 125 0 2 0 
2 126 1 125  
2 127 1 125  
1 128 0 3 0 
2 129 1 128  
2 130 1 128  
2 131 1 128  
1 132 0 4 0 
2 133 1 132  
2 134 1 132  
2 135 1 132  
2 136 1 132  
1 137 0 5 0 
2 138 1 137  
2 139 1 137  
2 140 1 137  
2 141 1 137  
2 142 1 137  
1 143 0 6 0 
2 144 1 143  
2 145 1 143  
2 146 1 143  
2 147 1 143  
2 148 1 143  
2 149 1 143  
1 150 0 8 0 
2 151 1 150  
2 152 1 150  
2 153 1 150  
2 154 1 150  
2 155 1 150  
2 156 1 150  
2 157 1 150  
2 158 1 150  
1 159 0 9 0 
2 160 1 159  
2 161 1 159  
2 162 1 159  
2 163 1 159  
2 164 1 159  
2 165 1 159  
2 166 1 159  
2 167 1 159  
2 168 1 159  
1 169 0 9 0 
2 170 1 169  
2 171 1 169  
2 172 1 169  
2 173 1 169  
2 174 1 169  
2 175 1 169  
2 176 1 169  
2 177 1 169  
2 178 1 169  
1 179 0 10 0 
2 180 1 179  
2 181 1 179  
2 182 1 179  
2 183 1 179  
2 184 1 179  
2 185 1 179  
2 186 1 179  
2 187 1 179  
2 188 1 179  
2 189 1 179  
1 190 0 9 0 
2 191 1 190  
2 192 1 190  
2 193 1 190  
2 194 1 190  
2 195 1 190  
2 196 1 190  
2 197 1 190  
2 198 1 190  
2 199 1 190  
1 200 0 12 0 
2 201 1 200  
2 202 1 200  
2 203 1 200  
2 204 1 200  
2 205 1 200  
2 206 1 200  
2 207 1 200  
2 208 1 200  
2 209 1 200  
2 210 1 200  
2 211 1 200  
2 212 1 200  
1 213 0 8 0 
2 214 1 213  
2 215 1 213  
2 216 1 213  
2 217 1 213  
2 218 1 213  
2 219 1 213  
2 220 1 213  
2 221 1 213  
1 222 0 1 0 
1 223 0 2 0 
2 224 1 223  
2 225 1 223  
1 226 0 5 0 
2 227 1 226  
2 228 1 226  
2 229 1 226  
2 230 1 226  
2 231 1 226  
1 232 0 5 0 
2 233 1 232  
2 234 1 232  
2 235 1 232  
2 236 1 232  
2 237 1 232  
1 238 0 5 0 
2 239 1 238  
2 240 1 238  
2 241 1 238  
2 242 1 238  
2 243 1 238  
1 244 0 5 0 
2 245 1 244  
2 246 1 244  
2 247 1 244  
2 248 1 244  
2 249 1 244  
1 250 0 6 0 
2 251 1 250  
2 252 1 250  
2 253 1 250  
2 254 1 250  
2 255 1 250  
2 256 1 250  
1 257 0 6 0 
2 258 1 257  
2 259 1 257  
2 260 1 257  
2 261 1 257  
2 262 1 257  
2 263 1 257  
1 264 0 5 0 
2 265 1 264  
2 266 1 264  
2 267 1 264  
2 268 1 264  
2 269 1 264  
1 270 0 3 0 
2 271 1 270  
2 272 1 270  
2 273 1 270  
1 274 0 8 0 
2 275 1 274  
2 276 1 274  
2 277 1 274  
2 278 1 274  
2 279 1 274  
2 280 1 274  
2 281 1 274  
2 282 1 274  
1 283 0 10 0 
2 284 1 283  
2 285 1 283  
2 286 1 283  
2 287 1 283  
2 288 1 283  
2 289 1 283  
2 290 1 283  
2 291 1 283  
2 292 1 283  
2 293 1 283  
1 294 0 8 0 
2 295 1 294  
2 296 1 294  
2 297 1 294  
2 298 1 294  
2 299 1 294  
2 300 1 294  
2 301 1 294  
2 302 1 294  
1 303 0 7 0 
2 304 1 303  
2 305 1 303  
2 306 1 303  
2 307 1 303  
2 308 1 303  
2 309 1 303  
2 310 1 303  
1 311 0 5 0 
2 312 1 311  
2 313 1 311  
2 314 1 311  
2 315 1 311  
2 316 1 311  
1 317 0 4 0 
2 318 1 317  
2 319 1 317  
2 320 1 317  
2 321 1 317  
1 322 0 3 0 
2 323 1 322  
2 324 1 322  
2 325 1 322  
1 326 0 2 0 
2 327 1 326  
2 328 1 326  
1 329 0 1 0 
1 330 0 12 0 
2 331 1 330  
2 332 1 330  
2 333 1 330  
2 334 1 330  
2 335 1 330  
2 336 1 330  
2 337 1 330  
2 338 1 330  
2 339 1 330  
2 340 1 330  
2 341 1 330  
2 342 1 330  
1 343 0 5 0 
2 344 1 343  
2 345 1 343  
2 346 1 343  
2 347 1 343  
2 348 1 343  
1 349 0 1 0 
1 350 0 2 0 
2 351 1 350  
2 352 1 350  
0 655 0 9 1 51 
2 656 1 655  
2 657 1 655  
2 658 1 655  
2 659 1 655  
2 660 1 655  
2 661 1 655  
2 662 1 655  
2 663 1 655  
2 664 1 655  
0 665 5 4 1 52 
2 666 1 665  
2 667 1 665  
2 668 1 665  
2 669 1 665  
0 670 0 8 1 59 
2 671 1 670  
2 672 1 670  
2 673 1 670  
2 674 1 670  
2 675 1 670  
2 676 1 670  
2 677 1 670  
2 678 1 670  
0 679 5 3 1 60 
2 680 1 679  
2 681 1 679  
2 682 1 679  
0 683 0 2 1 69 
2 684 1 683  
2 685 1 683  
0 686 5 3 1 70 
2 687 1 686  
2 688 1 686  
2 689 1 686  
0 690 0 8 1 71 
2 691 1 690  
2 692 1 690  
2 693 1 690  
2 694 1 690  
2 695 1 690  
2 696 1 690  
2 697 1 690  
2 698 1 690  
0 699 0 2 1 78 
2 700 1 699  
2 701 1 699  
0 702 5 3 1 79 
2 703 1 702  
2 704 1 702  
2 705 1 702  
0 706 0 8 1 80 
2 707 1 706  
2 708 1 706  
2 709 1 706  
2 710 1 706  
2 711 1 706  
2 712 1 706  
2 713 1 706  
2 714 1 706  
0 715 0 8 1 88 
2 716 1 715  
2 717 1 715  
2 718 1 715  
2 719 1 715  
2 720 1 715  
2 721 1 715  
2 722 1 715  
2 723 1 715  
0 724 5 2 1 89 
2 725 1 724  
2 726 1 724  
0 727 0 8 1 98 
2 728 1 727  
2 729 1 727  
2 730 1 727  
2 731 1 727  
2 732 1 727  
2 733 1 727  
2 734 1 727  
2 735 1 727  
0 736 5 3 1 99 
2 737 1 736  
2 738 1 736  
2 739 1 736  
0 740 0 8 1 108 
2 741 1 740  
2 742 1 740  
2 743 1 740  
2 744 1 740  
2 745 1 740  
2 746 1 740  
2 747 1 740  
2 748 1 740  
0 749 5 3 1 109 
2 750 1 749  
2 751 1 749  
2 752 1 749  
0 753 0 9 1 117 
2 754 1 753  
2 755 1 753  
2 756 1 753  
2 757 1 753  
2 758 1 753  
2 759 1 753  
2 760 1 753  
2 761 1 753  
2 762 1 753  
0 763 5 4 1 118 
2 764 1 763  
2 765 1 763  
2 766 1 763  
2 767 1 763  
0 768 3 1 2 258 265 
0 769 5 2 1 2 
2 770 1 769  
2 771 1 769  
0 772 0 6 1 3 
2 773 1 772  
2 774 1 772  
2 775 1 772  
2 776 1 772  
2 777 1 772  
2 778 1 772  
0 779 5 2 1 4 
2 780 1 779  
2 781 1 779  
0 782 0 3 1 14 
2 783 1 782  
2 784 1 782  
2 785 1 782  
0 786 5 6 1 15 
2 787 1 786  
2 788 1 786  
2 789 1 786  
2 790 1 786  
2 791 1 786  
2 792 1 786  
0 793 7 1 2 16 21 
0 794 5 3 1 22 
2 795 1 794  
2 796 1 794  
2 797 1 794  
0 798 0 4 1 23 
2 799 1 798  
2 800 1 798  
2 801 1 798  
2 802 1 798  
0 803 5 16 1 24 
2 804 1 803  
2 805 1 803  
2 806 1 803  
2 807 1 803  
2 808 1 803  
2 809 1 803  
2 810 1 803  
2 811 1 803  
2 812 1 803  
2 813 1 803  
2 814 1 803  
2 815 1 803  
2 816 1 803  
2 817 1 803  
2 818 1 803  
2 819 1 803  
0 820 5 1 1 34 
0 821 0 3 1 35 
2 822 1 821  
2 823 1 821  
2 824 1 821  
0 825 5 3 1 36 
2 826 1 825  
2 827 1 825  
2 828 1 825  
0 829 7 2 2 37 42 
2 830 1 829  
2 831 1 829  
0 832 5 2 1 43 
2 833 1 832  
2 834 1 832  
0 835 3 1 2 44 46 
0 836 0 2 1 47 
2 837 1 836  
2 838 1 836  
0 839 5 2 1 48 
2 840 1 839  
2 841 1 839  
0 842 5 2 1 53 
2 843 1 842  
2 844 1 842  
0 845 0 2 1 61 
2 846 1 845  
2 847 1 845  
0 848 5 2 1 62 
2 849 1 848  
2 850 1 848  
0 851 0 2 1 72 
2 852 1 851  
2 853 1 851  
0 854 5 3 1 73 
2 855 1 854  
2 856 1 854  
2 857 1 854  
0 858 0 2 1 90 
2 859 1 858  
2 860 1 858  
0 861 5 2 1 91 
2 862 1 861  
2 863 1 861  
0 864 0 2 1 100 
2 865 1 864  
2 866 1 864  
0 867 5 2 1 101 
2 868 1 867  
2 869 1 867  
0 870 5 3 1 110 
2 871 1 870  
2 872 1 870  
2 873 1 870  
0 874 0 2 1 5 
2 875 1 874  
2 876 1 874  
0 877 0 2 1 74 
2 878 1 877  
2 879 1 877  
0 880 0 2 1 111 
2 881 1 880  
2 882 1 880  
0 883 5 2 1 25 
2 884 1 883  
2 885 1 883  
0 886 0 2 1 191 
2 887 1 886  
2 888 1 886  
0 889 5 1 1 201 
0 890 7 1 2 26 202 
0 891 6 1 2 27 203 
0 892 7 2 2 28 180 
2 893 1 892  
2 894 1 892  
0 895 5 1 1 29 
0 896 3 16 2 349 38 
2 897 1 896  
2 898 1 896  
2 899 1 896  
2 900 1 896  
2 901 1 896  
2 902 1 896  
2 903 1 896  
2 904 1 896  
2 905 1 896  
2 906 1 896  
2 907 1 896  
2 908 1 896  
2 909 1 896  
2 910 1 896  
2 911 1 896  
2 912 1 896  
0 913 6 1 2 6 17 
0 914 6 1 3 7 30 39 
0 915 5 1 1 31 
0 916 5 1 1 40 
0 917 0 2 1 181 
2 918 1 917  
2 919 1 917  
0 920 5 2 1 214 
2 921 1 920  
2 922 1 920  
0 923 0 2 1 344 
2 924 1 923  
2 925 1 923  
0 926 0 2 1 227 
2 927 1 926  
2 928 1 926  
0 929 0 2 1 233 
2 930 1 929  
2 931 1 929  
0 932 0 2 1 239 
2 933 1 932  
2 934 1 932  
0 935 0 2 1 245 
2 936 1 935  
2 937 1 935  
0 938 0 2 1 251 
2 939 1 938  
2 940 1 938  
0 941 0 2 1 259 
2 942 1 941  
2 943 1 941  
0 944 0 2 1 266 
2 945 1 944  
2 946 1 944  
0 947 0 2 1 271 
2 948 1 947  
2 949 1 947  
0 950 0 2 1 54 
2 951 1 950  
2 952 1 950  
0 953 0 2 1 63 
2 954 1 953  
2 955 1 953  
0 956 0 2 1 64 
2 957 1 956  
2 958 1 956  
0 959 0 2 1 102 
2 960 1 959  
2 961 1 959  
0 962 0 2 1 103 
2 963 1 962  
2 964 1 962  
0 965 0 2 1 331 
2 966 1 965  
2 967 1 965  
0 1067 7 1 2 252 768 
0 1117 3 16 2 820 32 
2 1118 1 1117  
2 1119 1 1117  
2 1120 1 1117  
2 1121 1 1117  
2 1122 1 1117  
2 1123 1 1117  
2 1124 1 1117  
2 1125 1 1117  
2 1126 1 1117  
2 1127 1 1117  
2 1128 1 1117  
2 1129 1 1117  
2 1130 1 1117  
2 1131 1 1117  
2 1132 1 1117  
2 1133 1 1117  
0 1179 3 1 2 895 170 
0 1196 5 1 1 793 
0 1197 3 4 2 915 8 
2 1198 1 1197  
2 1199 1 1197  
2 1200 1 1197  
2 1201 1 1197  
0 1202 7 16 2 913 914 
2 1203 1 1202  
2 1204 1 1202  
2 1205 1 1202  
2 1206 1 1202  
2 1207 1 1202  
2 1208 1 1202  
2 1209 1 1202  
2 1210 1 1202  
2 1211 1 1202  
2 1212 1 1202  
2 1213 1 1202  
2 1214 1 1202  
2 1215 1 1202  
2 1216 1 1202  
2 1217 1 1202  
2 1218 1 1202  
0 1219 3 4 2 916 9 
2 1220 1 1219  
2 1221 1 1219  
2 1222 1 1219  
2 1223 1 1219  
0 1250 7 1 3 843 849 855 
0 1251 6 1 2 228 656 
0 1252 6 1 2 234 671 
0 1253 6 1 2 240 691 
0 1254 6 1 2 246 707 
0 1255 6 1 2 253 716 
0 1256 6 1 2 260 728 
0 1257 6 1 2 267 741 
0 1258 6 1 2 272 754 
0 1259 5 1 1 927 
0 1260 5 1 1 930 
0 1261 5 1 1 933 
0 1262 5 1 1 936 
0 1263 6 1 2 680 687 
0 1264 6 2 2 737 750 
2 1265 1 1264  
2 1266 1 1264  
0 1267 6 1 2 684 700 
0 1268 0 2 1 666 
2 1269 1 1268  
2 1270 1 1268  
0 1271 5 1 1 954 
0 1272 5 1 1 960 
0 1273 0 2 1 840 
2 1274 1 1273  
2 1275 1 1273  
0 1276 0 2 1 841 
2 1277 1 1276  
2 1278 1 1276  
0 1279 0 2 1 783 
2 1280 1 1279  
2 1281 1 1279  
0 1298 0 3 1 826 
2 1299 1 1298  
2 1300 1 1298  
2 1301 1 1298  
0 1302 0 3 1 833 
2 1303 1 1302  
2 1304 1 1302  
2 1305 1 1302  
0 1306 7 8 2 780 835 
2 1307 1 1306  
2 1308 1 1306  
2 1309 1 1306  
2 1310 1 1306  
2 1311 1 1306  
2 1312 1 1306  
2 1313 1 1306  
2 1314 1 1306  
0 1315 7 6 3 781 837 834 
2 1316 1 1315  
2 1317 1 1315  
2 1318 1 1315  
2 1319 1 1315  
2 1320 1 1315  
2 1321 1 1315  
0 1322 7 2 2 770 838 
2 1323 1 1322  
2 1324 1 1322  
0 1325 7 2 3 773 787 799 
2 1326 1 1325  
2 1327 1 1325  
0 1328 6 2 3 774 788 800 
2 1329 1 1328  
2 1330 1 1328  
0 1331 6 2 2 775 789 
2 1332 1 1331  
2 1333 1 1331  
0 1334 0 2 1 875 
2 1335 1 1334  
2 1336 1 1334  
0 1337 6 1 3 784 795 49 
0 1338 6 1 3 844 850 856 
0 1339 5 1 1 957 
0 1340 7 2 3 862 868 871 
2 1341 1 1340  
2 1342 1 1340  
0 1343 6 1 3 863 869 872 
0 1344 5 1 1 963 
0 1345 5 1 1 804 
0 1346 5 1 1 805 
0 1347 5 1 1 806 
0 1348 5 1 1 807 
0 1349 5 1 1 808 
0 1350 5 1 1 809 
0 1351 5 1 1 810 
0 1352 5 1 1 811 
0 1353 3 4 2 884 887 
2 1354 1 1353  
2 1355 1 1353  
2 1356 1 1353  
2 1357 1 1353  
0 1358 4 4 2 885 888 
2 1359 1 1358  
2 1360 1 1358  
2 1361 1 1358  
2 1362 1 1358  
0 1363 0 2 1 893 
2 1364 1 1363  
2 1365 1 1363  
0 1366 5 2 1 894 
2 1367 1 1366  
2 1368 1 1366  
0 1369 0 14 1 822 
2 1370 1 1369  
2 1371 1 1369  
2 1372 1 1369  
2 1373 1 1369  
2 1374 1 1369  
2 1375 1 1369  
2 1376 1 1369  
2 1377 1 1369  
2 1378 1 1369  
2 1379 1 1369  
2 1380 1 1369  
2 1381 1 1369  
2 1382 1 1369  
2 1383 1 1369  
0 1384 0 16 1 827 
2 1385 1 1384  
2 1386 1 1384  
2 1387 1 1384  
2 1388 1 1384  
2 1389 1 1384  
2 1390 1 1384  
2 1391 1 1384  
2 1392 1 1384  
2 1393 1 1384  
2 1394 1 1384  
2 1395 1 1384  
2 1396 1 1384  
2 1397 1 1384  
2 1398 1 1384  
2 1399 1 1384  
2 1400 1 1384  
0 1401 5 1 1 897 
0 1402 5 1 1 898 
0 1403 5 1 1 899 
0 1404 5 1 1 900 
0 1405 5 1 1 901 
0 1406 5 1 1 902 
0 1407 5 1 1 903 
0 1408 5 1 1 904 
0 1409 3 16 2 10 1196 
2 1410 1 1409  
2 1411 1 1409  
2 1412 1 1409  
2 1413 1 1409  
2 1414 1 1409  
2 1415 1 1409  
2 1416 1 1409  
2 1417 1 1409  
2 1418 1 1409  
2 1419 1 1409  
2 1420 1 1409  
2 1421 1 1409  
2 1422 1 1409  
2 1423 1 1409  
2 1424 1 1409  
2 1425 1 1409  
0 1426 5 1 1 830 
0 1427 5 1 1 831 
0 1452 7 6 3 771 785 796 
2 1453 1 1452  
2 1454 1 1452  
2 1455 1 1452  
2 1456 1 1452  
2 1457 1 1452  
2 1458 1 1452  
0 1459 5 1 1 918 
0 1460 5 1 1 966 
0 1461 3 2 2 921 924 
2 1462 1 1461  
2 1463 1 1461  
0 1464 4 2 2 922 925 
2 1465 1 1464  
2 1466 1 1464  
0 1467 5 1 1 939 
0 1468 5 1 1 942 
0 1469 5 1 1 945 
0 1470 5 1 1 948 
0 1471 0 2 1 681 
2 1472 1 1471  
2 1473 1 1471  
0 1474 5 1 1 951 
0 1475 0 2 1 688 
2 1476 1 1475  
2 1477 1 1475  
0 1478 0 2 1 703 
2 1479 1 1478  
2 1480 1 1478  
0 1481 0 2 1 725 
2 1482 1 1481  
2 1483 1 1481  
0 1484 0 2 1 738 
2 1485 1 1484  
2 1486 1 1484  
0 1487 0 2 1 751 
2 1488 1 1487  
2 1489 1 1487  
0 1490 0 2 1 764 
2 1491 1 1490  
2 1492 1 1490  
0 1493 0 2 1 878 
2 1494 1 1493  
2 1495 1 1493  
0 1496 0 2 1 879 
2 1497 1 1496  
2 1498 1 1496  
0 1499 0 2 1 881 
2 1500 1 1499  
2 1501 1 1499  
0 1502 0 2 1 882 
2 1503 1 1502  
2 1504 1 1502  
0 1505 6 1 2 704 1250 
0 1507 7 1 4 1251 1252 1253 1254 
0 1508 7 1 4 1255 1256 1257 1258 
0 1509 6 1 2 931 1259 
0 1510 6 1 2 928 1260 
0 1511 6 1 2 937 1261 
0 1512 6 1 2 934 1262 
0 1520 7 3 2 657 1263 
2 1521 1 1520  
2 1522 1 1520  
2 1523 1 1520  
0 1562 7 16 2 876 1337 
2 1563 1 1562  
2 1564 1 1562  
2 1565 1 1562  
2 1566 1 1562  
2 1567 1 1562  
2 1568 1 1562  
2 1569 1 1562  
2 1570 1 1562  
2 1571 1 1562  
2 1572 1 1562  
2 1573 1 1562  
2 1574 1 1562  
2 1575 1 1562  
2 1576 1 1562  
2 1577 1 1562  
2 1578 1 1562  
0 1579 5 1 1 1118 
0 1580 7 1 2 812 1119 
0 1581 7 1 2 1338 1345 
0 1582 5 1 1 1120 
0 1583 7 1 2 813 1121 
0 1584 5 1 1 1122 
0 1585 7 1 2 814 1123 
0 1586 7 1 2 857 1347 
0 1587 5 1 1 1124 
0 1588 7 1 2 815 1125 
0 1589 7 1 2 81 1348 
0 1590 5 1 1 1126 
0 1591 7 1 2 816 1127 
0 1592 7 1 2 1343 1349 
0 1593 5 1 1 1128 
0 1594 7 1 2 817 1129 
0 1595 5 1 1 1130 
0 1596 7 1 2 818 1131 
0 1597 7 1 2 873 1351 
0 1598 5 1 1 1132 
0 1599 7 1 2 819 1133 
0 1600 7 1 2 119 1352 
0 1643 7 1 2 222 1401 
0 1644 7 1 2 224 1402 
0 1645 7 1 2 229 1403 
0 1646 7 1 2 235 1404 
0 1647 7 1 2 241 1405 
0 1648 7 1 2 247 1406 
0 1649 7 1 2 254 1407 
0 1650 7 1 2 261 1408 
0 1667 7 2 3 11 18 1426 
2 1668 1 1667  
2 1669 1 1667  
0 1670 7 2 3 12 19 1427 
2 1671 1 1670  
2 1672 1 1670  
0 1673 5 1 1 1203 
0 1674 5 1 1 1204 
0 1675 5 1 1 1205 
0 1676 5 1 1 1206 
0 1677 5 1 1 1207 
0 1678 5 1 1 1208 
0 1679 5 1 1 1209 
0 1680 5 1 1 1210 
0 1691 6 1 2 943 1467 
0 1692 6 1 2 940 1468 
0 1693 6 1 2 949 1469 
0 1694 6 1 2 946 1470 
3 1713 5 0 1 1505 
0 1714 7 1 2 92 1265 
0 1715 6 2 2 1509 1510 
2 1716 1 1715  
2 1717 1 1715  
0 1718 6 2 2 1511 1512 
2 1719 1 1718  
2 1720 1 1718  
0 1721 6 1 2 1507 1508 
0 1722 7 2 2 765 1341 
2 1723 1 1722  
2 1724 1 1722  
0 1725 6 1 2 766 1342 
0 1726 5 1 1 1269 
0 1727 6 1 2 1494 1271 
0 1728 5 1 1 1495 
0 1729 7 1 2 685 1270 
0 1730 6 1 2 1500 1272 
0 1731 5 1 1 1501 
0 1735 6 1 2 93 1266 
0 1736 5 1 1 1274 
0 1737 5 1 1 1277 
0 1738 6 8 2 1326 823 
2 1739 1 1738  
2 1740 1 1738  
2 1741 1 1738  
2 1742 1 1738  
2 1743 1 1738  
2 1744 1 1738  
2 1745 1 1738  
2 1746 1 1738  
0 1747 6 8 2 1327 828 
2 1748 1 1747  
2 1749 1 1747  
2 1750 1 1747  
2 1751 1 1747  
2 1752 1 1747  
2 1753 1 1747  
2 1754 1 1747  
2 1755 1 1747  
0 1756 6 4 3 776 1280 801 
2 1757 1 1756  
2 1758 1 1756  
2 1759 1 1756  
2 1760 1 1756  
0 1761 6 2 4 777 790 802 1303 
2 1762 1 1761  
2 1763 1 1761  
0 1764 6 1 2 1497 1339 
0 1765 5 1 1 1498 
0 1766 6 1 2 1503 1344 
0 1767 5 1 1 1504 
0 1768 5 1 1 1329 
0 1769 5 1 1 1335 
0 1770 5 1 1 1332 
0 1787 7 1 2 846 1579 
0 1788 7 1 2 151 1580 
0 1789 7 1 2 852 1582 
0 1790 7 1 2 160 1583 
0 1791 7 1 2 82 1584 
0 1792 7 1 2 55 1585 
0 1793 7 1 2 859 1587 
0 1794 7 1 2 847 1588 
0 1795 7 1 2 865 1590 
0 1796 7 1 2 853 1591 
0 1797 7 1 2 112 1593 
0 1798 7 1 2 83 1594 
0 1799 7 1 2 120 1595 
0 1800 7 1 2 860 1596 
0 1801 7 1 2 284 1598 
0 1802 7 1 2 866 1599 
0 1803 7 2 2 204 1364 
2 1804 1 1803  
2 1805 1 1803  
0 1806 7 2 2 889 1365 
2 1807 1 1806  
2 1808 1 1806  
0 1809 7 2 2 890 1367 
2 1810 1 1809  
2 1811 1 1809  
0 1812 7 2 2 891 1368 
2 1813 1 1812  
2 1814 1 1812  
0 1815 6 2 2 1299 1304 
2 1816 1 1815  
2 1817 1 1815  
0 1818 6 2 2 824 1305 
2 1819 1 1818  
2 1820 1 1818  
0 1821 6 2 3 778 1281 1179 
2 1822 1 1821  
2 1823 1 1821  
0 1824 6 8 3 791 797 1300 
2 1825 1 1824  
2 1826 1 1824  
2 1827 1 1824  
2 1828 1 1824  
2 1829 1 1824  
2 1830 1 1824  
2 1831 1 1824  
2 1832 1 1824  
0 1833 6 8 2 792 1301 
2 1834 1 1833  
2 1835 1 1833  
2 1836 1 1833  
2 1837 1 1833  
2 1838 1 1833  
2 1839 1 1833  
2 1840 1 1833  
2 1841 1 1833  
0 1842 5 1 1 1370 
0 1843 5 1 1 1371 
0 1844 5 1 1 1372 
0 1845 5 1 1 1373 
0 1846 5 1 1 1374 
0 1847 5 1 1 1375 
0 1848 5 1 1 1376 
0 1849 5 1 1 1385 
0 1850 7 1 2 1386 905 
0 1851 5 1 1 1387 
0 1852 7 1 2 1388 906 
0 1853 5 1 1 1389 
0 1854 7 1 2 1390 907 
0 1855 5 1 1 1391 
0 1856 7 1 2 1392 908 
0 1857 5 1 1 1393 
0 1858 7 1 2 1394 909 
0 1859 5 1 1 1395 
0 1860 7 1 2 1396 910 
0 1861 5 1 1 1397 
0 1862 7 1 2 1398 911 
0 1863 5 1 1 1399 
0 1864 7 1 2 1400 912 
0 1869 7 1 2 1211 1410 
0 1870 4 2 2 56 1411 
2 1871 1 1870  
2 1872 1 1870  
0 1873 5 1 1 1307 
0 1874 7 1 2 1212 1412 
0 1875 4 2 2 65 1413 
2 1876 1 1875  
2 1877 1 1875  
0 1878 5 1 1 1308 
0 1879 7 1 2 1213 1414 
0 1880 4 2 2 75 1415 
2 1881 1 1880  
2 1882 1 1880  
0 1883 5 1 1 1309 
0 1884 7 1 2 1214 1416 
0 1885 4 2 2 84 1417 
2 1886 1 1885  
2 1887 1 1885  
0 1888 5 1 1 1310 
0 1889 7 1 2 1215 1418 
0 1890 4 2 2 94 1419 
2 1891 1 1890  
2 1892 1 1890  
0 1893 5 1 1 1323 
0 1894 7 1 2 1216 1420 
0 1895 4 2 2 104 1421 
2 1896 1 1895  
2 1897 1 1895  
0 1898 5 1 1 1316 
0 1899 7 1 2 1217 1422 
0 1900 4 2 2 113 1423 
2 1901 1 1900  
2 1902 1 1900  
0 1903 5 1 1 1317 
0 1904 7 1 2 1218 1424 
0 1905 4 2 2 121 1425 
2 1906 1 1905  
2 1907 1 1905  
0 1908 5 1 1 1318 
0 1909 7 2 2 1453 215 
2 1910 1 1909  
2 1911 1 1909  
0 1912 6 1 2 1454 216 
0 1913 7 3 3 1455 217 345 
2 1914 1 1913  
2 1915 1 1913  
2 1916 1 1913  
0 1917 6 4 3 1456 218 346 
2 1918 1 1917  
2 1919 1 1917  
2 1920 1 1917  
2 1921 1 1917  
0 1922 7 3 3 1457 219 347 
2 1923 1 1922  
2 1924 1 1922  
2 1925 1 1922  
0 1926 6 3 3 1458 220 348 
2 1927 1 1926  
2 1928 1 1926  
2 1929 1 1926  
0 1930 0 2 1 1465 
2 1931 1 1930  
2 1932 1 1930  
0 1933 6 2 2 1691 1692 
2 1934 1 1933  
2 1935 1 1933  
0 1936 6 2 2 1693 1694 
2 1937 1 1936  
2 1938 1 1936  
0 1939 5 1 1 1472 
0 1940 6 1 2 1473 1474 
0 1941 5 1 1 1476 
0 1942 5 1 1 1479 
0 1943 5 1 1 1482 
0 1944 5 1 1 1485 
0 1945 5 1 1 1488 
0 1946 5 1 1 1491 
3 1947 5 0 1 1714 
0 1960 6 1 2 955 1728 
0 1961 6 1 2 961 1731 
0 1966 7 1 2 1521 1278 
0 1981 6 1 2 958 1765 
0 1982 6 1 2 964 1767 
0 1983 7 2 2 1067 1768 
2 1984 1 1983  
2 1985 1 1983  
0 1986 3 1 3 1581 1787 1788 
0 1987 3 1 3 1586 1791 1792 
0 1988 3 1 3 1589 1793 1794 
0 1989 3 1 3 1592 1795 1796 
0 1990 3 1 3 1597 1799 1800 
0 1991 3 1 3 1600 1801 1802 
0 2022 7 1 2 85 1849 
0 2023 7 1 2 225 1850 
0 2024 7 1 2 95 1851 
0 2025 7 1 2 230 1852 
0 2026 7 1 2 105 1853 
0 2027 7 1 2 236 1854 
0 2028 7 1 2 114 1855 
0 2029 7 1 2 242 1856 
0 2030 7 1 2 122 1857 
0 2031 7 1 2 248 1858 
0 2032 7 1 2 285 1859 
0 2033 7 1 2 255 1860 
0 2034 7 1 2 295 1861 
0 2035 7 1 2 262 1862 
0 2036 7 1 2 304 1863 
0 2037 7 1 2 268 1864 
0 2038 0 4 1 1668 
2 2039 1 2038  
2 2040 1 2038  
2 2041 1 2038  
2 2042 1 2038  
0 2043 5 8 1 1669 
2 2044 1 2043  
2 2045 1 2043  
2 2046 1 2043  
2 2047 1 2043  
2 2048 1 2043  
2 2049 1 2043  
2 2050 1 2043  
2 2051 1 2043  
0 2052 0 4 1 1671 
2 2053 1 2052  
2 2054 1 2052  
2 2055 1 2052  
2 2056 1 2052  
0 2057 5 8 1 1672 
2 2058 1 2057  
2 2059 1 2057  
2 2060 1 2057  
2 2061 1 2057  
2 2062 1 2057  
2 2063 1 2057  
2 2064 1 2057  
2 2065 1 2057  
0 2068 7 2 3 57 1198 1869 
2 2069 1 2068  
2 2070 1 2068  
0 2073 7 2 3 66 1199 1874 
2 2074 1 2073  
2 2075 1 2073  
0 2078 7 2 3 76 1200 1879 
2 2079 1 2078  
2 2080 1 2078  
0 2083 7 2 3 86 1201 1884 
2 2084 1 2083  
2 2085 1 2083  
0 2088 7 2 3 96 1220 1889 
2 2089 1 2088  
2 2090 1 2088  
0 2093 7 2 3 106 1221 1894 
2 2094 1 2093  
2 2095 1 2093  
0 2098 7 2 3 115 1222 1899 
2 2099 1 2098  
2 2100 1 2098  
0 2103 7 2 3 123 1223 1904 
2 2104 1 2103  
2 2105 1 2103  
0 2121 5 1 1 1563 
0 2122 5 1 1 1564 
0 2123 5 1 1 1565 
0 2124 5 1 1 1566 
0 2125 5 1 1 1567 
0 2126 5 1 1 1568 
0 2127 5 1 1 1569 
0 2128 5 1 1 1570 
0 2133 6 1 2 952 1939 
0 2134 6 1 2 1480 1941 
0 2135 6 1 2 1477 1942 
0 2136 6 1 2 1486 1943 
0 2137 6 1 2 1483 1944 
0 2138 6 1 2 1492 1945 
0 2139 6 1 2 1489 1946 
0 2141 5 1 1 1934 
0 2142 5 1 1 1937 
0 2143 5 1 1 1739 
0 2144 7 1 2 1740 1748 
0 2145 5 1 1 1749 
0 2146 6 1 2 1727 1960 
0 2147 6 1 2 1730 1961 
0 2148 7 1 4 1723 1267 667 67 
0 2149 5 1 1 1741 
0 2150 7 1 2 1742 1750 
0 2151 5 1 1 1751 
0 2152 5 1 1 1743 
0 2153 5 1 1 1752 
0 2154 7 1 2 1744 1753 
0 2155 5 1 1 1745 
0 2156 5 1 1 1754 
0 2157 7 1 2 1746 1755 
0 2158 0 16 1 1762 
2 2159 1 2158  
2 2160 1 2158  
2 2161 1 2158  
2 2162 1 2158  
2 2163 1 2158  
2 2164 1 2158  
2 2165 1 2158  
2 2166 1 2158  
2 2167 1 2158  
2 2168 1 2158  
2 2169 1 2158  
2 2170 1 2158  
2 2171 1 2158  
2 2172 1 2158  
2 2173 1 2158  
2 2174 1 2158  
0 2175 0 2 1 1763 
2 2176 1 2175  
2 2177 1 2175  
0 2178 6 1 2 1764 1981 
0 2179 6 1 2 1766 1982 
0 2180 5 1 1 1757 
0 2181 7 1 2 1758 1330 
0 2183 5 1 1 1759 
0 2184 7 1 2 1333 1760 
0 2185 6 2 2 1359 1813 
2 2186 1 2185  
2 2187 1 2185  
0 2188 6 2 2 1360 1810 
2 2189 1 2188  
2 2190 1 2188  
0 2191 6 2 2 1354 1814 
2 2192 1 2191  
2 2193 1 2191  
0 2194 6 2 2 1355 1811 
2 2195 1 2194  
2 2196 1 2194  
0 2197 6 2 2 1361 1807 
2 2198 1 2197  
2 2199 1 2197  
0 2200 6 2 2 1362 1804 
2 2201 1 2200  
2 2202 1 2200  
0 2203 6 2 2 1356 1808 
2 2204 1 2203  
2 2205 1 2203  
0 2206 6 2 2 1357 1805 
2 2207 1 2206  
2 2208 1 2206  
0 2209 5 1 1 1816 
0 2210 5 1 1 1819 
0 2211 7 1 2 1817 1820 
0 2212 0 8 1 1822 
2 2213 1 2212  
2 2214 1 2212  
2 2215 1 2212  
2 2216 1 2212  
2 2217 1 2212  
2 2218 1 2212  
2 2219 1 2212  
2 2220 1 2212  
0 2221 0 8 1 1823 
2 2222 1 2221  
2 2223 1 2221  
2 2224 1 2221  
2 2225 1 2221  
2 2226 1 2221  
2 2227 1 2221  
2 2228 1 2221  
2 2229 1 2221  
0 2230 5 1 1 1834 
0 2231 5 1 1 1835 
0 2232 5 1 1 1836 
0 2233 5 1 1 1837 
0 2234 5 1 1 1825 
0 2235 5 1 1 1826 
0 2236 5 1 1 1827 
0 2237 5 1 1 1828 
0 2238 3 1 3 2022 1643 2023 
0 2239 3 1 3 2024 1644 2025 
0 2240 3 1 3 2026 1645 2027 
0 2241 3 1 3 2028 1646 2029 
0 2242 3 1 3 2030 1647 2031 
0 2243 3 1 3 2032 1648 2033 
0 2244 3 1 3 2034 1649 2035 
0 2245 3 1 3 2036 1650 2037 
0 2270 7 2 2 1986 1673 
2 2271 1 2270  
2 2272 1 2270  
0 2277 7 2 2 1987 1675 
2 2278 1 2277  
2 2279 1 2277  
0 2282 7 2 2 1988 1676 
2 2283 1 2282  
2 2284 1 2282  
0 2287 7 2 2 1989 1677 
2 2288 1 2287  
2 2289 1 2287  
0 2294 7 2 2 1990 1679 
2 2295 1 2294  
2 2296 1 2294  
0 2299 7 2 2 1991 1680 
2 2300 1 2299  
2 2301 1 2299  
0 2304 0 2 1 1918 
2 2305 1 2304  
2 2306 1 2304  
0 2307 7 2 2 1931 351 
2 2308 1 2307  
2 2309 1 2307  
0 2310 6 2 2 1932 352 
2 2311 1 2310  
2 2312 1 2310  
0 2313 0 2 1 1716 
2 2314 1 2313  
2 2315 1 2313  
0 2316 0 2 1 1719 
2 2317 1 2316  
2 2318 1 2316  
0 2319 0 2 1 1717 
2 2320 1 2319  
2 2321 1 2319  
0 2322 0 2 1 1720 
2 2323 1 2322  
2 2324 1 2322  
0 2325 6 2 2 1940 2133 
2 2326 1 2325  
2 2327 1 2325  
0 2328 6 2 2 2134 2135 
2 2329 1 2328  
2 2330 1 2328  
0 2331 6 2 2 2136 2137 
2 2332 1 2331  
2 2333 1 2331  
0 2334 6 2 2 2138 2139 
2 2335 1 2334  
2 2336 1 2334  
0 2341 6 1 2 1938 2141 
0 2342 6 1 2 1935 2142 
0 2347 7 1 2 726 2144 
0 2348 7 1 3 2146 701 1726 
0 2349 7 1 2 755 2147 
0 2350 7 1 2 2148 1275 
0 2351 7 1 2 739 2150 
0 2352 7 1 2 1735 2153 
0 2353 7 1 2 767 2154 
0 2354 7 1 2 1725 2156 
0 2355 7 1 2 752 2157 
0 2374 5 1 1 2178 
0 2375 5 1 1 2179 
0 2376 7 2 2 1522 2180 
2 2377 1 2376  
2 2378 1 2376  
0 2379 7 2 2 1721 2181 
2 2380 1 2379  
2 2381 1 2379  
0 2398 7 1 2 668 2211 
0 2417 7 1 3 2058 231 1873 
0 2418 7 1 3 2059 275 1311 
0 2419 7 1 2 2053 2238 
0 2420 7 1 3 2060 237 1878 
0 2421 7 1 3 2061 276 1312 
0 2422 7 1 2 2054 2239 
0 2425 7 1 3 2062 243 1883 
0 2426 7 1 3 2063 277 1313 
0 2427 7 1 2 2055 2240 
0 2430 7 1 3 2064 249 1888 
0 2431 7 1 3 2065 278 1314 
0 2432 7 1 2 2056 2241 
0 2435 7 1 3 2044 256 1893 
0 2436 7 1 3 2045 279 1324 
0 2437 7 1 2 2039 2242 
0 2438 7 1 3 2046 263 1898 
0 2439 7 1 3 2047 280 1319 
0 2440 7 1 2 2040 2243 
0 2443 7 1 3 2048 269 1903 
0 2444 7 1 3 2049 281 1320 
0 2445 7 1 2 2041 2244 
0 2448 7 1 3 2050 273 1908 
0 2449 7 1 3 2051 282 1321 
0 2450 7 1 2 2042 2245 
0 2467 5 1 1 2314 
0 2468 5 1 1 2317 
0 2469 5 1 1 2320 
0 2470 5 1 1 2323 
0 2471 6 2 2 2341 2342 
2 2472 1 2471  
2 2473 1 2471  
0 2474 5 1 1 2326 
0 2475 5 1 1 2329 
0 2476 5 1 1 2332 
0 2477 5 1 1 2335 
0 2478 3 1 2 2348 1729 
0 2481 5 1 1 2176 
0 2482 7 1 2 2177 1336 
0 2483 7 2 2 2349 2183 
2 2484 1 2483  
2 2485 1 2483  
0 2486 7 1 2 2374 1346 
0 2487 7 1 2 2375 1350 
0 2488 0 8 1 2186 
2 2489 1 2488  
2 2490 1 2488  
2 2491 1 2488  
2 2492 1 2488  
2 2493 1 2488  
2 2494 1 2488  
2 2495 1 2488  
2 2496 1 2488  
0 2497 0 8 1 2189 
2 2498 1 2497  
2 2499 1 2497  
2 2500 1 2497  
2 2501 1 2497  
2 2502 1 2497  
2 2503 1 2497  
2 2504 1 2497  
2 2505 1 2497  
0 2506 0 8 1 2192 
2 2507 1 2506  
2 2508 1 2506  
2 2509 1 2506  
2 2510 1 2506  
2 2511 1 2506  
2 2512 1 2506  
2 2513 1 2506  
2 2514 1 2506  
0 2515 0 8 1 2195 
2 2516 1 2515  
2 2517 1 2515  
2 2518 1 2515  
2 2519 1 2515  
2 2520 1 2515  
2 2521 1 2515  
2 2522 1 2515  
2 2523 1 2515  
0 2524 0 8 1 2198 
2 2525 1 2524  
2 2526 1 2524  
2 2527 1 2524  
2 2528 1 2524  
2 2529 1 2524  
2 2530 1 2524  
2 2531 1 2524  
2 2532 1 2524  
0 2533 0 8 1 2201 
2 2534 1 2533  
2 2535 1 2533  
2 2536 1 2533  
2 2537 1 2533  
2 2538 1 2533  
2 2539 1 2533  
2 2540 1 2533  
2 2541 1 2533  
0 2542 0 8 1 2204 
2 2543 1 2542  
2 2544 1 2542  
2 2545 1 2542  
2 2546 1 2542  
2 2547 1 2542  
2 2548 1 2542  
2 2549 1 2542  
2 2550 1 2542  
0 2551 0 8 1 2207 
2 2552 1 2551  
2 2553 1 2551  
2 2554 1 2551  
2 2555 1 2551  
2 2556 1 2551  
2 2557 1 2551  
2 2558 1 2551  
2 2559 1 2551  
0 2560 0 8 1 2187 
2 2561 1 2560  
2 2562 1 2560  
2 2563 1 2560  
2 2564 1 2560  
2 2565 1 2560  
2 2566 1 2560  
2 2567 1 2560  
2 2568 1 2560  
0 2569 0 8 1 2190 
2 2570 1 2569  
2 2571 1 2569  
2 2572 1 2569  
2 2573 1 2569  
2 2574 1 2569  
2 2575 1 2569  
2 2576 1 2569  
2 2577 1 2569  
0 2578 0 8 1 2193 
2 2579 1 2578  
2 2580 1 2578  
2 2581 1 2578  
2 2582 1 2578  
2 2583 1 2578  
2 2584 1 2578  
2 2585 1 2578  
2 2586 1 2578  
0 2587 0 8 1 2196 
2 2588 1 2587  
2 2589 1 2587  
2 2590 1 2587  
2 2591 1 2587  
2 2592 1 2587  
2 2593 1 2587  
2 2594 1 2587  
2 2595 1 2587  
0 2596 0 8 1 2199 
2 2597 1 2596  
2 2598 1 2596  
2 2599 1 2596  
2 2600 1 2596  
2 2601 1 2596  
2 2602 1 2596  
2 2603 1 2596  
2 2604 1 2596  
0 2605 0 8 1 2202 
2 2606 1 2605  
2 2607 1 2605  
2 2608 1 2605  
2 2609 1 2605  
2 2610 1 2605  
2 2611 1 2605  
2 2612 1 2605  
2 2613 1 2605  
0 2614 0 8 1 2205 
2 2615 1 2614  
2 2616 1 2614  
2 2617 1 2614  
2 2618 1 2614  
2 2619 1 2614  
2 2620 1 2614  
2 2621 1 2614  
2 2622 1 2614  
0 2623 0 8 1 2208 
2 2624 1 2623  
2 2625 1 2623  
2 2626 1 2623  
2 2627 1 2623  
2 2628 1 2623  
2 2629 1 2623  
2 2630 1 2623  
2 2631 1 2623  
0 2632 5 1 1 2213 
0 2633 7 1 2 2214 1838 
0 2634 5 1 1 2215 
0 2635 7 1 2 2216 1839 
0 2636 5 1 1 2217 
0 2637 7 1 2 2218 1840 
0 2638 5 1 1 2219 
0 2639 7 1 2 2220 1841 
0 2640 5 1 1 2222 
0 2641 7 1 2 2223 1829 
0 2642 5 1 1 2224 
0 2643 7 1 2 2225 1830 
0 2644 5 1 1 2226 
0 2645 7 1 2 2227 1831 
0 2646 5 1 1 2228 
0 2647 7 1 2 2229 1832 
0 2648 3 3 3 2271 1871 2069 
2 2649 1 2648  
2 2650 1 2648  
2 2651 1 2648  
0 2652 4 3 3 2272 1872 2070 
2 2653 1 2652  
2 2654 1 2652  
2 2655 1 2652  
0 2656 3 2 3 2417 2418 2419 
2 2657 1 2656  
2 2658 1 2656  
0 2659 3 2 3 2420 2421 2422 
2 2660 1 2659  
2 2661 1 2659  
0 2662 3 3 3 2278 1881 2079 
2 2663 1 2662  
2 2664 1 2662  
2 2665 1 2662  
0 2666 4 3 3 2279 1882 2080 
2 2667 1 2666  
2 2668 1 2666  
2 2669 1 2666  
0 2670 3 2 3 2425 2426 2427 
2 2671 1 2670  
2 2672 1 2670  
0 2673 3 3 3 2283 1886 2084 
2 2674 1 2673  
2 2675 1 2673  
2 2676 1 2673  
0 2677 4 3 3 2284 1887 2085 
2 2678 1 2677  
2 2679 1 2677  
2 2680 1 2677  
0 2681 3 2 3 2430 2431 2432 
2 2682 1 2681  
2 2683 1 2681  
0 2684 3 3 3 2288 1891 2089 
2 2685 1 2684  
2 2686 1 2684  
2 2687 1 2684  
0 2688 4 3 3 2289 1892 2090 
2 2689 1 2688  
2 2690 1 2688  
2 2691 1 2688  
0 2692 3 4 3 2435 2436 2437 
2 2693 1 2692  
2 2694 1 2692  
2 2695 1 2692  
2 2696 1 2692  
0 2697 3 4 3 2438 2439 2440 
2 2698 1 2697  
2 2699 1 2697  
2 2700 1 2697  
2 2701 1 2697  
0 2702 3 3 3 2295 1901 2099 
2 2703 1 2702  
2 2704 1 2702  
2 2705 1 2702  
0 2706 4 3 3 2296 1902 2100 
2 2707 1 2706  
2 2708 1 2706  
2 2709 1 2706  
0 2710 3 4 3 2443 2444 2445 
2 2711 1 2710  
2 2712 1 2710  
2 2713 1 2710  
2 2714 1 2710  
0 2715 3 3 3 2300 1906 2104 
2 2716 1 2715  
2 2717 1 2715  
2 2718 1 2715  
0 2719 4 3 3 2301 1907 2105 
2 2720 1 2719  
2 2721 1 2719  
2 2722 1 2719  
0 2723 3 4 3 2448 2449 2450 
2 2724 1 2723  
2 2725 1 2723  
2 2726 1 2723  
2 2727 1 2723  
0 2728 5 1 1 2305 
0 2729 5 1 1 2159 
0 2730 7 1 2 1571 2160 
0 2731 5 1 1 2161 
0 2732 7 1 2 1572 2162 
0 2733 5 1 1 2163 
0 2734 7 1 2 1573 2164 
0 2735 5 1 1 2165 
0 2736 7 1 2 1574 2166 
0 2737 5 1 1 2167 
0 2738 7 1 2 1575 2168 
0 2739 5 1 1 2169 
0 2740 7 1 2 1576 2170 
0 2741 5 1 1 2171 
0 2742 7 1 2 1577 2172 
0 2743 5 1 1 2173 
0 2744 7 1 2 1578 2174 
0 2745 3 1 3 2377 1984 2380 
0 2746 4 1 3 2378 1985 2381 
0 2748 6 1 2 2318 2467 
0 2749 6 1 2 2315 2468 
0 2750 6 1 2 2324 2469 
0 2751 6 1 2 2321 2470 
0 2754 6 1 2 2330 2474 
0 2755 6 1 2 2327 2475 
0 2756 6 1 2 2336 2476 
0 2757 6 1 2 2333 2477 
0 2758 7 2 2 1523 2481 
2 2759 1 2758  
2 2760 1 2758  
0 2761 7 2 2 1724 2482 
2 2762 1 2761  
2 2763 1 2761  
0 2764 7 2 2 2478 1770 
2 2765 1 2764  
2 2766 1 2764  
0 2768 3 1 3 2486 1789 1790 
0 2769 3 1 3 2487 1797 1798 
0 2898 7 1 2 669 2633 
0 2899 7 1 2 682 2635 
0 2900 7 1 2 689 2637 
0 2901 7 1 2 705 2639 
0 2962 5 1 1 2746 
0 2966 6 1 2 2748 2749 
0 2967 6 2 2 2750 2751 
2 2968 1 2967  
2 2969 1 2967  
0 2970 0 2 1 2472 
2 2971 1 2970  
2 2972 1 2970  
0 2973 6 3 2 2754 2755 
2 2974 1 2973  
2 2975 1 2973  
2 2976 1 2973  
0 2977 6 2 2 2756 2757 
2 2978 1 2977  
2 2979 1 2977  
0 2980 7 1 2 2473 2143 
0 2984 5 1 1 2489 
0 2985 5 1 1 2498 
0 2986 5 1 1 2507 
0 2987 5 1 1 2516 
0 2988 5 1 1 2525 
0 2989 5 1 1 2534 
0 2990 5 1 1 2543 
0 2991 5 1 1 2552 
0 2992 5 1 1 2490 
0 2993 5 1 1 2499 
0 2994 5 1 1 2508 
0 2995 5 1 1 2517 
0 2996 5 1 1 2526 
0 2997 5 1 1 2535 
0 2998 5 1 1 2544 
0 2999 5 1 1 2553 
0 3000 5 1 1 2491 
0 3001 5 1 1 2500 
0 3002 5 1 1 2509 
0 3003 5 1 1 2518 
0 3004 5 1 1 2527 
0 3005 5 1 1 2536 
0 3006 5 1 1 2545 
0 3007 5 1 1 2554 
0 3008 5 1 1 2492 
0 3009 5 1 1 2501 
0 3010 5 1 1 2510 
0 3011 5 1 1 2519 
0 3012 5 1 1 2528 
0 3013 5 1 1 2537 
0 3014 5 1 1 2546 
0 3015 5 1 1 2555 
0 3016 5 1 1 2493 
0 3017 5 1 1 2502 
0 3018 5 1 1 2511 
0 3019 5 1 1 2520 
0 3020 5 1 1 2529 
0 3021 5 1 1 2538 
0 3022 5 1 1 2547 
0 3023 5 1 1 2556 
0 3024 5 1 1 2494 
0 3025 5 1 1 2503 
0 3026 5 1 1 2512 
0 3027 5 1 1 2521 
0 3028 5 1 1 2530 
0 3029 5 1 1 2539 
0 3030 5 1 1 2548 
0 3031 5 1 1 2557 
0 3032 5 1 1 2495 
0 3033 5 1 1 2504 
0 3034 5 1 1 2513 
0 3035 5 1 1 2522 
0 3036 5 1 1 2531 
0 3037 5 1 1 2540 
0 3038 5 1 1 2549 
0 3039 5 1 1 2558 
0 3040 5 1 1 2496 
0 3041 5 1 1 2505 
0 3042 5 1 1 2514 
0 3043 5 1 1 2523 
0 3044 5 1 1 2532 
0 3045 5 1 1 2541 
0 3046 5 1 1 2550 
0 3047 5 1 1 2559 
0 3048 5 1 1 2561 
0 3049 5 1 1 2570 
0 3050 5 1 1 2579 
0 3051 5 1 1 2588 
0 3052 5 1 1 2597 
0 3053 5 1 1 2606 
0 3054 5 1 1 2615 
0 3055 5 1 1 2624 
0 3056 5 1 1 2562 
0 3057 5 1 1 2571 
0 3058 5 1 1 2580 
0 3059 5 1 1 2589 
0 3060 5 1 1 2598 
0 3061 5 1 1 2607 
0 3062 5 1 1 2616 
0 3063 5 1 1 2625 
0 3064 5 1 1 2563 
0 3065 5 1 1 2572 
0 3066 5 1 1 2581 
0 3067 5 1 1 2590 
0 3068 5 1 1 2599 
0 3069 5 1 1 2608 
0 3070 5 1 1 2617 
0 3071 5 1 1 2626 
0 3072 5 1 1 2564 
0 3073 5 1 1 2573 
0 3074 5 1 1 2582 
0 3075 5 1 1 2591 
0 3076 5 1 1 2600 
0 3077 5 1 1 2609 
0 3078 5 1 1 2618 
0 3079 5 1 1 2627 
0 3080 5 1 1 2565 
0 3081 5 1 1 2574 
0 3082 5 1 1 2583 
0 3083 5 1 1 2592 
0 3084 5 1 1 2601 
0 3085 5 1 1 2610 
0 3086 5 1 1 2619 
0 3087 5 1 1 2628 
0 3088 5 1 1 2566 
0 3089 5 1 1 2575 
0 3090 5 1 1 2584 
0 3091 5 1 1 2593 
0 3092 5 1 1 2602 
0 3093 5 1 1 2611 
0 3094 5 1 1 2620 
0 3095 5 1 1 2629 
0 3096 5 1 1 2567 
0 3097 5 1 1 2576 
0 3098 5 1 1 2585 
0 3099 5 1 1 2594 
0 3100 5 1 1 2603 
0 3101 5 1 1 2612 
0 3102 5 1 1 2621 
0 3103 5 1 1 2630 
0 3104 5 1 1 2568 
0 3105 5 1 1 2577 
0 3106 5 1 1 2586 
0 3107 5 1 1 2595 
0 3108 5 1 1 2604 
0 3109 5 1 1 2613 
0 3110 5 1 1 2622 
0 3111 5 1 1 2631 
0 3112 0 2 1 2657 
2 3113 1 3112  
2 3114 1 3112  
0 3115 5 2 1 2658 
2 3116 1 3115  
2 3117 1 3115  
0 3118 5 1 1 2653 
0 3119 7 2 2 2768 1674 
2 3120 1 3119  
2 3121 1 3119  
0 3122 0 2 1 2660 
2 3123 1 3122  
2 3124 1 3122  
0 3125 5 2 1 2661 
2 3126 1 3125  
2 3127 1 3125  
0 3128 0 2 1 2671 
2 3129 1 3128  
2 3130 1 3128  
0 3131 5 2 1 2672 
2 3132 1 3131  
2 3133 1 3131  
0 3134 5 1 1 2667 
0 3135 0 2 1 2682 
2 3136 1 3135  
2 3137 1 3135  
0 3138 5 2 1 2683 
2 3139 1 3138  
2 3140 1 3138  
0 3141 5 1 1 2678 
0 3142 0 2 1 2693 
2 3143 1 3142  
2 3144 1 3142  
0 3145 5 2 1 2694 
2 3146 1 3145  
2 3147 1 3145  
0 3148 5 1 1 2689 
0 3149 7 2 2 2769 1678 
2 3150 1 3149  
2 3151 1 3149  
0 3152 0 2 1 2698 
2 3153 1 3152  
2 3154 1 3152  
0 3155 5 2 1 2699 
2 3156 1 3155  
2 3157 1 3155  
0 3158 0 2 1 2711 
2 3159 1 3158  
2 3160 1 3158  
0 3161 5 2 1 2712 
2 3162 1 3161  
2 3163 1 3161  
0 3164 5 1 1 2707 
0 3165 0 2 1 2724 
2 3166 1 3165  
2 3167 1 3165  
0 3168 5 2 1 2725 
2 3169 1 3168  
2 3170 1 3168  
0 3171 5 1 1 2720 
0 3172 7 2 2 1910 2649 
2 3173 1 3172  
2 3174 1 3172  
0 3175 7 2 2 1914 2663 
2 3176 1 3175  
2 3177 1 3175  
0 3178 7 2 2 1915 2674 
2 3179 1 3178  
2 3180 1 3178  
0 3181 7 2 2 1916 2685 
2 3182 1 3181  
2 3183 1 3181  
0 3184 7 2 2 1923 2703 
2 3185 1 3184  
2 3186 1 3184  
0 3187 7 2 2 1924 2716 
2 3188 1 3187  
2 3189 1 3187  
0 3190 5 1 1 2695 
0 3191 5 1 1 2700 
0 3192 5 1 1 2713 
0 3193 5 1 1 2726 
0 3194 7 1 5 2696 2701 2714 2727 1459 
3 3195 6 0 2 2745 2962 
0 3196 5 1 1 2966 
0 3206 3 1 3 2980 2145 2347 
0 3207 7 1 2 124 2984 
0 3208 7 1 2 161 2985 
0 3209 7 1 2 152 2986 
0 3210 7 1 2 144 2987 
0 3211 7 1 2 138 2988 
0 3212 7 1 2 133 2989 
0 3213 7 1 2 129 2990 
0 3214 7 1 2 126 2991 
0 3215 7 1 2 127 2992 
0 3216 7 1 2 658 2993 
0 3217 7 1 2 162 2994 
0 3218 7 1 2 153 2995 
0 3219 7 1 2 145 2996 
0 3220 7 1 2 139 2997 
0 3221 7 1 2 134 2998 
0 3222 7 1 2 130 2999 
0 3223 7 1 2 131 3000 
0 3224 7 1 2 672 3001 
0 3225 7 1 2 659 3002 
0 3226 7 1 2 163 3003 
0 3227 7 1 2 154 3004 
0 3228 7 1 2 146 3005 
0 3229 7 1 2 140 3006 
0 3230 7 1 2 135 3007 
0 3231 7 1 2 136 3008 
0 3232 7 1 2 692 3009 
0 3233 7 1 2 673 3010 
0 3234 7 1 2 660 3011 
0 3235 7 1 2 164 3012 
0 3236 7 1 2 155 3013 
0 3237 7 1 2 147 3014 
0 3238 7 1 2 141 3015 
0 3239 7 1 2 142 3016 
0 3240 7 1 2 708 3017 
0 3241 7 1 2 693 3018 
0 3242 7 1 2 674 3019 
0 3243 7 1 2 661 3020 
0 3244 7 1 2 165 3021 
0 3245 7 1 2 156 3022 
0 3246 7 1 2 148 3023 
0 3247 7 1 2 149 3024 
0 3248 7 1 2 717 3025 
0 3249 7 1 2 709 3026 
0 3250 7 1 2 694 3027 
0 3251 7 1 2 675 3028 
0 3252 7 1 2 662 3029 
0 3253 7 1 2 166 3030 
0 3254 7 1 2 157 3031 
0 3255 7 1 2 158 3032 
0 3256 7 1 2 729 3033 
0 3257 7 1 2 718 3034 
0 3258 7 1 2 710 3035 
0 3259 7 1 2 695 3036 
0 3260 7 1 2 676 3037 
0 3261 7 1 2 663 3038 
0 3262 7 1 2 167 3039 
0 3263 7 1 2 168 3040 
0 3264 7 1 2 742 3041 
0 3265 7 1 2 730 3042 
0 3266 7 1 2 719 3043 
0 3267 7 1 2 711 3044 
0 3268 7 1 2 696 3045 
0 3269 7 1 2 677 3046 
0 3270 7 1 2 664 3047 
0 3271 7 1 2 286 3048 
0 3272 7 1 2 678 3049 
0 3273 7 1 2 697 3050 
0 3274 7 1 2 712 3051 
0 3275 7 1 2 720 3052 
0 3276 7 1 2 731 3053 
0 3277 7 1 2 743 3054 
0 3278 7 1 2 756 3055 
0 3279 7 1 2 296 3056 
0 3280 7 1 2 698 3057 
0 3281 7 1 2 713 3058 
0 3282 7 1 2 721 3059 
0 3283 7 1 2 732 3060 
0 3284 7 1 2 744 3061 
0 3285 7 1 2 757 3062 
0 3286 7 1 2 287 3063 
0 3287 7 1 2 305 3064 
0 3288 7 1 2 714 3065 
0 3289 7 1 2 722 3066 
0 3290 7 1 2 733 3067 
0 3291 7 1 2 745 3068 
0 3292 7 1 2 758 3069 
0 3293 7 1 2 288 3070 
0 3294 7 1 2 297 3071 
0 3295 7 1 2 312 3072 
0 3296 7 1 2 723 3073 
0 3297 7 1 2 734 3074 
0 3298 7 1 2 746 3075 
0 3299 7 1 2 759 3076 
0 3300 7 1 2 289 3077 
0 3301 7 1 2 298 3078 
0 3302 7 1 2 306 3079 
0 3303 7 1 2 318 3080 
0 3304 7 1 2 735 3081 
0 3305 7 1 2 747 3082 
0 3306 7 1 2 760 3083 
0 3307 7 1 2 290 3084 
0 3308 7 1 2 299 3085 
0 3309 7 1 2 307 3086 
0 3310 7 1 2 313 3087 
0 3311 7 1 2 323 3088 
0 3312 7 1 2 748 3089 
0 3313 7 1 2 761 3090 
0 3314 7 1 2 291 3091 
0 3315 7 1 2 300 3092 
0 3316 7 1 2 308 3093 
0 3317 7 1 2 314 3094 
0 3318 7 1 2 319 3095 
0 3319 7 1 2 327 3096 
0 3320 7 1 2 762 3097 
0 3321 7 1 2 292 3098 
0 3322 7 1 2 301 3099 
0 3323 7 1 2 309 3100 
0 3324 7 1 2 315 3101 
0 3325 7 1 2 320 3102 
0 3326 7 1 2 324 3103 
0 3327 7 1 2 329 3104 
0 3328 7 1 2 293 3105 
0 3329 7 1 2 302 3106 
0 3330 7 1 2 310 3107 
0 3331 7 1 2 316 3108 
0 3332 7 1 2 321 3109 
0 3333 7 1 2 325 3110 
0 3334 7 1 2 328 3111 
0 3383 7 1 5 3190 3191 3192 3193 919 
0 3384 0 2 1 2978 
2 3385 1 3384  
2 3386 1 3384  
0 3387 7 1 2 3196 1736 
0 3388 7 1 2 2979 2149 
0 3389 7 1 2 2974 1737 
0 3390 4 1 8 3207 3208 3209 3210 3211 3212 3213 3214 
0 3391 4 1 8 3215 3216 3217 3218 3219 3220 3221 3222 
0 3392 4 1 8 3223 3224 3225 3226 3227 3228 3229 3230 
0 3393 4 1 8 3231 3232 3233 3234 3235 3236 3237 3238 
0 3394 4 1 8 3239 3240 3241 3242 3243 3244 3245 3246 
0 3395 4 1 8 3247 3248 3249 3250 3251 3252 3253 3254 
0 3396 4 1 8 3255 3256 3257 3258 3259 3260 3261 3262 
0 3397 4 1 8 3263 3264 3265 3266 3267 3268 3269 3270 
0 3398 4 1 8 3271 3272 3273 3274 3275 3276 3277 3278 
0 3399 4 1 8 3279 3280 3281 3282 3283 3284 3285 3286 
0 3400 4 1 8 3287 3288 3289 3290 3291 3292 3293 3294 
0 3401 4 1 8 3295 3296 3297 3298 3299 3300 3301 3302 
0 3402 4 1 8 3303 3304 3305 3306 3307 3308 3309 3310 
0 3403 4 1 8 3311 3312 3313 3314 3315 3316 3317 3318 
0 3404 4 1 8 3319 3320 3321 3322 3323 3324 3325 3326 
0 3405 4 1 8 3327 3328 3329 3330 3331 3332 3333 3334 
0 3406 7 1 2 3206 2641 
0 3407 7 2 3 171 2650 3113 
2 3408 1 3407  
2 3409 1 3407  
0 3410 7 2 3 182 2651 3116 
2 3411 1 3410  
2 3412 1 3410  
0 3413 7 1 3 192 2654 3117 
0 3414 7 1 3 205 2655 3114 
0 3415 3 3 3 3120 1876 2074 
2 3416 1 3415  
2 3417 1 3415  
2 3418 1 3415  
0 3419 4 3 3 3121 1877 2075 
2 3420 1 3419  
2 3421 1 3419  
2 3422 1 3419  
0 3423 7 2 3 172 2664 3129 
2 3424 1 3423  
2 3425 1 3423  
0 3426 7 2 3 183 2665 3132 
2 3427 1 3426  
2 3428 1 3426  
0 3429 7 1 3 193 2668 3133 
0 3430 7 1 3 206 2669 3130 
0 3431 7 2 3 173 2675 3136 
2 3432 1 3431  
2 3433 1 3431  
0 3434 7 2 3 184 2676 3139 
2 3435 1 3434  
2 3436 1 3434  
0 3437 7 1 3 194 2679 3140 
0 3438 7 1 3 207 2680 3137 
0 3439 7 2 3 174 2686 3143 
2 3440 1 3439  
2 3441 1 3439  
0 3442 7 2 3 185 2687 3146 
2 3443 1 3442  
2 3444 1 3442  
0 3445 7 1 3 195 2690 3147 
0 3446 7 1 3 208 2691 3144 
0 3447 3 3 3 3150 1896 2094 
2 3448 1 3447  
2 3449 1 3447  
2 3450 1 3447  
0 3451 4 3 3 3151 1897 2095 
2 3452 1 3451  
2 3453 1 3451  
2 3454 1 3451  
0 3455 7 2 3 175 2704 3159 
2 3456 1 3455  
2 3457 1 3455  
0 3458 7 2 3 186 2705 3162 
2 3459 1 3458  
2 3460 1 3458  
0 3461 7 1 3 196 2708 3163 
0 3462 7 1 3 209 2709 3160 
0 3463 7 2 3 176 2717 3166 
2 3464 1 3463  
2 3465 1 3463  
0 3466 7 2 3 187 2718 3169 
2 3467 1 3466  
2 3468 1 3466  
0 3469 7 1 3 197 2721 3170 
0 3470 7 1 3 210 2722 3167 
0 3471 3 1 2 3194 3383 
0 3472 0 2 1 2968 
2 3473 1 3472  
2 3474 1 3472  
0 3475 0 2 1 2971 
2 3476 1 3475  
2 3477 1 3475  
0 3478 0 2 1 2969 
2 3479 1 3478  
2 3480 1 3478  
0 3481 0 2 1 2972 
2 3482 1 3481  
2 3483 1 3481  
0 3484 0 2 1 2975 
2 3485 1 3484  
2 3486 1 3484  
0 3487 0 2 1 2976 
2 3488 1 3487  
2 3489 1 3487  
0 3490 0 2 1 3173 
2 3491 1 3490  
2 3492 1 3490  
0 3493 0 2 1 3174 
2 3494 1 3493  
2 3495 1 3493  
0 3496 0 2 1 3176 
2 3497 1 3496  
2 3498 1 3496  
0 3499 0 2 1 3177 
2 3500 1 3499  
2 3501 1 3499  
0 3502 0 2 1 3179 
2 3503 1 3502  
2 3504 1 3502  
0 3505 0 2 1 3180 
2 3506 1 3505  
2 3507 1 3505  
0 3508 0 2 1 3182 
2 3509 1 3508  
2 3510 1 3508  
0 3511 0 2 1 3183 
2 3512 1 3511  
2 3513 1 3511  
0 3514 0 2 1 3185 
2 3515 1 3514  
2 3516 1 3514  
0 3517 0 2 1 3186 
2 3518 1 3517  
2 3519 1 3517  
0 3520 0 2 1 3188 
2 3521 1 3520  
2 3522 1 3520  
0 3523 0 2 1 3189 
2 3524 1 3523  
2 3525 1 3523  
0 3534 4 1 2 3387 2350 
0 3535 3 1 3 3388 2151 2351 
0 3536 4 1 2 3389 1966 
0 3537 7 1 2 3390 2209 
0 3538 7 1 2 3398 2210 
0 3539 7 1 2 3391 1842 
0 3540 7 1 2 3399 1377 
0 3541 7 1 2 3392 1843 
0 3542 7 1 2 3400 1378 
0 3543 7 1 2 3393 1844 
0 3544 7 1 2 3401 1379 
0 3545 7 1 2 3394 1845 
0 3546 7 1 2 3402 1380 
0 3547 7 1 2 3395 1846 
0 3548 7 1 2 3403 1381 
0 3549 7 1 2 3396 1847 
0 3550 7 1 2 3404 1382 
0 3551 7 1 2 3397 1848 
0 3552 7 1 2 3405 1383 
0 3557 3 1 3 3413 3414 3118 
0 3568 3 1 3 3429 3430 3134 
0 3573 3 1 3 3437 3438 3141 
0 3578 3 1 3 3445 3446 3148 
0 3589 3 1 3 3461 3462 3164 
0 3594 3 1 3 3469 3470 3171 
0 3605 7 1 2 3471 2728 
0 3626 5 1 1 3479 
0 3627 5 1 1 3482 
0 3628 5 1 1 3488 
0 3629 5 1 1 3485 
0 3630 5 1 1 3473 
0 3631 5 1 1 3476 
0 3632 7 1 2 3536 2152 
0 3633 7 1 2 3534 2155 
0 3634 3 1 3 3537 3538 2398 
0 3635 3 1 2 3539 3540 
0 3636 3 1 2 3541 3542 
0 3637 3 1 2 3543 3544 
0 3638 3 1 2 3545 3546 
0 3639 3 1 2 3547 3548 
0 3640 3 1 2 3549 3550 
0 3641 3 1 2 3551 3552 
0 3642 7 1 2 3535 2643 
0 3643 3 1 2 3408 3411 
0 3644 4 1 2 3409 3412 
0 3645 7 2 3 177 3416 3123 
2 3646 1 3645  
2 3647 1 3645  
0 3648 7 2 3 188 3417 3126 
2 3649 1 3648  
2 3650 1 3648  
0 3651 7 1 3 198 3420 3127 
0 3652 7 1 3 211 3421 3124 
0 3653 5 1 1 3422 
0 3654 3 2 2 3424 3427 
2 3655 1 3654  
2 3656 1 3654  
0 3657 4 1 2 3425 3428 
0 3658 3 2 2 3432 3435 
2 3659 1 3658  
2 3660 1 3658  
0 3661 4 1 2 3433 3436 
0 3662 3 1 2 3440 3443 
0 3663 4 1 2 3441 3444 
0 3664 7 2 3 178 3448 3153 
2 3665 1 3664  
2 3666 1 3664  
0 3667 7 2 3 189 3449 3156 
2 3668 1 3667  
2 3669 1 3667  
0 3670 7 1 3 199 3452 3157 
0 3671 7 1 3 212 3453 3154 
0 3672 5 1 1 3454 
0 3673 3 2 2 3456 3459 
2 3674 1 3673  
2 3675 1 3673  
0 3676 4 1 2 3457 3460 
0 3677 3 2 2 3464 3467 
2 3678 1 3677  
2 3679 1 3677  
0 3680 4 1 2 3465 3468 
0 3681 5 1 1 3494 
0 3682 7 2 2 1911 3418 
2 3683 1 3682  
2 3684 1 3682  
0 3685 5 1 1 3497 
0 3686 5 1 1 3500 
0 3687 5 1 1 3503 
0 3688 5 1 1 3506 
0 3689 5 1 1 3512 
0 3690 7 2 2 1925 3450 
2 3691 1 3690  
2 3692 1 3690  
0 3693 5 1 1 3518 
0 3694 5 1 1 3521 
0 3695 5 1 1 3524 
0 3696 5 1 1 3515 
0 3697 0 2 1 3385 
2 3698 1 3697  
2 3699 1 3697  
0 3700 0 2 1 3386 
2 3701 1 3700  
2 3702 1 3700  
0 3703 5 1 1 3491 
0 3704 5 1 1 3509 
0 3705 6 1 2 3477 3630 
0 3706 6 1 2 3474 3631 
0 3707 6 1 2 3483 3626 
0 3708 6 1 2 3480 3627 
0 3711 3 1 3 3632 2352 2353 
0 3712 3 1 3 3633 2354 2355 
0 3713 7 1 2 3634 2632 
0 3714 7 1 2 3635 2634 
0 3715 7 1 2 3636 2636 
0 3716 7 1 2 3637 2638 
0 3717 7 1 2 3638 2640 
0 3718 7 1 2 3639 2642 
0 3719 7 1 2 3640 2644 
0 3720 7 1 2 3641 2646 
0 3721 7 5 2 3644 3557 
2 3722 1 3721  
2 3723 1 3721  
2 3724 1 3721  
2 3725 1 3721  
2 3726 1 3721  
0 3731 3 1 3 3651 3652 3653 
0 3734 7 3 2 3657 3568 
2 3735 1 3734  
2 3736 1 3734  
2 3737 1 3734  
0 3740 7 2 2 3661 3573 
2 3741 1 3740  
2 3742 1 3740  
0 3743 7 5 2 3663 3578 
2 3744 1 3743  
2 3745 1 3743  
2 3746 1 3743  
2 3747 1 3743  
2 3748 1 3743  
0 3753 3 1 3 3670 3671 3672 
0 3756 7 3 2 3676 3589 
2 3757 1 3756  
2 3758 1 3756  
2 3759 1 3756  
0 3762 7 2 2 3680 3594 
2 3763 1 3762  
2 3764 1 3762  
0 3765 5 1 1 3643 
0 3766 5 1 1 3662 
0 3773 6 1 2 3705 3706 
0 3774 6 1 2 3707 3708 
0 3775 6 1 2 3701 3628 
0 3776 5 1 1 3702 
0 3777 6 1 2 3698 3629 
0 3778 5 1 1 3699 
0 3779 7 1 2 3712 2645 
0 3780 7 1 2 3711 2647 
0 3786 3 2 2 3646 3649 
2 3787 1 3786  
2 3788 1 3786  
0 3789 4 1 2 3647 3650 
0 3800 3 2 2 3665 3668 
2 3801 1 3800  
2 3802 1 3800  
0 3803 4 1 2 3666 3669 
0 3809 7 2 2 3655 1919 
2 3810 1 3809  
2 3811 1 3809  
0 3812 7 2 2 3659 1920 
2 3813 1 3812  
2 3814 1 3812  
0 3815 7 2 2 3674 1927 
2 3816 1 3815  
2 3817 1 3815  
0 3818 7 2 2 3678 1928 
2 3819 1 3818  
2 3820 1 3818  
0 3821 0 2 1 3683 
2 3822 1 3821  
2 3823 1 3821  
0 3824 0 2 1 3684 
2 3825 1 3824  
2 3826 1 3824  
0 3827 0 2 1 3691 
2 3828 1 3827  
2 3829 1 3827  
0 3830 0 2 1 3692 
2 3831 1 3830  
2 3832 1 3830  
3 3833 6 0 2 3773 3774 
0 3834 6 1 2 3489 3776 
0 3835 6 1 2 3486 3778 
0 3838 7 4 2 3789 3731 
2 3839 1 3838  
2 3840 1 3838  
2 3841 1 3838  
2 3842 1 3838  
0 3845 7 4 2 3803 3753 
2 3846 1 3845  
2 3847 1 3845  
2 3848 1 3845  
2 3849 1 3845  
0 3850 0 2 1 3722 
2 3851 1 3850  
2 3852 1 3850  
0 3855 0 2 1 3735 
2 3856 1 3855  
2 3857 1 3855  
0 3858 0 2 1 3741 
2 3859 1 3858  
2 3860 1 3858  
0 3861 0 2 1 3744 
2 3862 1 3861  
2 3863 1 3861  
0 3865 0 2 1 3757 
2 3866 1 3865  
2 3867 1 3865  
0 3868 0 2 1 3763 
2 3869 1 3868  
2 3870 1 3868  
0 3884 6 1 2 3775 3834 
0 3885 6 1 2 3777 3835 
0 3894 6 1 2 3723 3787 
0 3895 6 1 2 3745 3801 
0 3898 5 1 1 3822 
0 3899 5 1 1 3825 
0 3906 5 1 1 3831 
0 3911 5 1 1 3828 
0 3912 7 1 2 3788 1912 
0 3913 0 2 1 3813 
2 3914 1 3913  
2 3915 1 3913  
0 3916 7 1 2 3802 1921 
0 3917 0 2 1 3819 
2 3918 1 3917  
2 3919 1 3917  
0 3920 5 1 1 3810 
0 3921 0 2 1 3820 
2 3922 1 3921  
2 3923 1 3921  
0 3924 5 1 1 3884 
0 3925 5 1 1 3885 
0 3926 7 3 4 3724 3839 3736 3742 
2 3927 1 3926  
2 3928 1 3926  
2 3929 1 3926  
0 3930 6 1 3 3725 3840 3656 
0 3931 6 1 4 3660 3841 3737 3726 
0 3932 7 2 4 3746 3846 3758 3764 
2 3933 1 3932  
2 3934 1 3932  
0 3935 6 1 3 3747 3847 3675 
0 3936 6 1 4 3679 3848 3759 3748 
0 3937 0 2 1 3842 
2 3938 1 3937  
2 3939 1 3937  
0 3940 0 2 1 3849 
2 3941 1 3940  
2 3942 1 3940  
0 3947 5 1 1 3912 
0 3948 5 1 1 3916 
0 3950 0 2 1 3851 
2 3951 1 3950  
2 3952 1 3950  
0 3953 0 2 1 3852 
2 3954 1 3953  
2 3955 1 3953  
0 3956 0 2 1 3856 
2 3957 1 3956  
2 3958 1 3956  
0 3959 0 2 1 3857 
2 3960 1 3959  
2 3961 1 3959  
0 3962 0 2 1 3859 
2 3963 1 3962  
2 3964 1 3962  
0 3965 0 2 1 3860 
2 3966 1 3965  
2 3967 1 3965  
0 3968 0 2 1 3862 
2 3969 1 3968  
2 3970 1 3968  
0 3971 0 2 1 3863 
2 3972 1 3971  
2 3973 1 3971  
0 3974 0 2 1 3866 
2 3975 1 3974  
2 3976 1 3974  
0 3977 0 2 1 3867 
2 3978 1 3977  
2 3979 1 3977  
0 3980 0 2 1 3869 
2 3981 1 3980  
2 3982 1 3980  
0 3983 0 2 1 3870 
2 3984 1 3983  
2 3985 1 3983  
3 3987 6 0 2 3924 3925 
0 3992 6 2 4 3765 3894 3930 3931 
2 3993 1 3992  
2 3994 1 3992  
0 3996 6 2 4 3766 3895 3935 3936 
2 3997 1 3996  
2 3998 1 3996  
0 4013 5 1 1 3922 
3 4028 7 0 2 3933 3927 
0 4029 6 1 2 3954 3681 
0 4030 6 1 2 3960 3686 
0 4031 6 1 2 3966 3688 
0 4032 6 1 2 3972 3689 
0 4033 6 1 2 3978 3693 
0 4034 6 1 2 3984 3695 
0 4035 0 2 1 3928 
2 4036 1 4035  
2 4037 1 4035  
0 4042 5 1 1 3955 
0 4043 5 1 1 3957 
0 4044 6 1 2 3958 3685 
0 4045 5 1 1 3961 
0 4046 5 1 1 3963 
0 4047 6 1 2 3964 3687 
0 4048 5 1 1 3967 
0 4049 5 1 1 3973 
0 4050 5 1 1 3979 
0 4051 5 1 1 3981 
0 4052 6 1 2 3982 3694 
0 4053 5 1 1 3985 
0 4054 5 1 1 3975 
0 4055 6 1 2 3976 3696 
0 4056 7 1 2 3934 2306 
0 4057 5 1 1 3951 
0 4058 6 1 2 3952 3703 
0 4059 0 2 1 3938 
2 4060 1 4059  
2 4061 1 4059  
0 4062 0 2 1 3939 
2 4063 1 4062  
2 4064 1 4062  
0 4065 5 1 1 3969 
0 4066 6 1 2 3970 3704 
0 4067 0 2 1 3941 
2 4068 1 4067  
2 4069 1 4067  
0 4070 0 2 1 3942 
2 4071 1 4070  
2 4072 1 4070  
0 4073 6 1 2 3929 3997 
0 4074 5 1 1 3993 
0 4075 6 1 2 3495 4042 
0 4076 6 1 2 3501 4045 
0 4077 6 1 2 3507 4048 
0 4078 6 1 2 3513 4049 
0 4079 6 1 2 3519 4050 
0 4080 6 1 2 3525 4053 
0 4085 6 1 2 3498 4043 
0 4086 6 1 2 3504 4046 
0 4088 6 1 2 3522 4051 
0 4090 6 1 2 3516 4054 
0 4091 7 2 2 3998 1929 
2 4092 1 4091  
2 4093 1 4091  
0 4094 3 3 2 3605 4056 
2 4095 1 4094  
2 4096 1 4094  
2 4097 1 4094  
0 4098 6 1 2 3492 4057 
0 4101 6 1 2 3510 4065 
0 4104 7 1 2 4073 4074 
0 4105 6 1 2 4075 4029 
0 4106 6 1 2 4063 3899 
0 4107 6 1 2 4076 4030 
0 4108 6 1 2 4077 4031 
0 4109 6 1 2 4078 4032 
0 4110 6 1 2 4071 3906 
0 4111 6 1 2 4079 4033 
0 4112 6 1 2 4080 4034 
0 4113 5 1 1 4060 
0 4114 6 1 2 4061 3898 
0 4115 5 1 1 4064 
0 4116 6 2 2 4085 4044 
2 4117 1 4116  
2 4118 1 4116  
0 4119 6 2 2 4086 4047 
2 4120 1 4119  
2 4121 1 4119  
0 4122 5 1 1 4072 
0 4123 6 2 2 4088 4052 
2 4124 1 4123  
2 4125 1 4123  
0 4126 5 1 1 4068 
0 4127 6 1 2 4069 3911 
0 4128 6 5 2 4090 4055 
2 4129 1 4128  
2 4130 1 4128  
2 4131 1 4128  
2 4132 1 4128  
2 4133 1 4128  
0 4139 6 2 2 4098 4058 
2 4140 1 4139  
2 4141 1 4139  
0 4142 6 2 2 4101 4066 
2 4143 1 4142  
2 4144 1 4142  
3 4145 5 0 1 4104 
0 4146 5 1 1 4105 
0 4147 6 1 2 3826 4115 
0 4148 5 1 1 4107 
0 4149 5 1 1 4108 
0 4150 5 1 1 4109 
0 4151 6 1 2 3832 4122 
0 4152 5 1 1 4111 
0 4153 5 1 1 4112 
0 4154 6 1 2 3823 4113 
0 4161 6 1 2 3829 4126 
0 4167 0 6 1 4092 
2 4168 1 4167  
2 4169 1 4167  
2 4170 1 4167  
2 4171 1 4167  
2 4172 1 4167  
2 4173 1 4167  
0 4174 0 4 1 4095 
2 4175 1 4174  
2 4176 1 4174  
2 4177 1 4174  
2 4178 1 4174  
0 4182 0 2 1 4093 
2 4183 1 4182  
2 4184 1 4182  
0 4186 7 2 2 332 4096 
2 4187 1 4186  
2 4188 1 4186  
0 4189 7 1 2 4146 2230 
0 4190 6 1 2 4147 4106 
0 4191 7 1 2 4148 2232 
0 4192 7 1 2 4149 2233 
0 4193 7 1 2 4150 2234 
0 4194 6 1 2 4151 4110 
0 4195 7 1 2 4152 2236 
0 4196 7 1 2 4153 2237 
0 4197 6 2 2 4154 4114 
2 4198 1 4197  
2 4199 1 4197  
0 4200 0 2 1 4117 
2 4201 1 4200  
2 4202 1 4200  
0 4203 0 5 1 4118 
2 4204 1 4203  
2 4205 1 4203  
2 4206 1 4203  
2 4207 1 4203  
2 4208 1 4203  
0 4209 0 3 1 4120 
2 4210 1 4209  
2 4211 1 4209  
2 4212 1 4209  
0 4213 0 4 1 4121 
2 4214 1 4213  
2 4215 1 4213  
2 4216 1 4213  
2 4217 1 4213  
0 4218 6 4 2 4161 4127 
2 4219 1 4218  
2 4220 1 4218  
2 4221 1 4218  
2 4222 1 4218  
0 4223 0 4 1 4124 
2 4224 1 4223  
2 4225 1 4223  
2 4226 1 4223  
2 4227 1 4223  
0 4238 7 1 2 4129 3918 
0 4239 5 1 1 4140 
0 4241 5 1 1 4143 
0 4242 7 2 2 333 4125 
2 4243 1 4242  
2 4244 1 4242  
0 4247 0 2 1 4130 
2 4248 1 4247  
2 4249 1 4247  
0 4251 4 1 3 3713 4189 2898 
0 4252 5 1 1 4190 
0 4253 4 1 3 3715 4191 2900 
0 4254 4 1 3 3716 4192 2901 
0 4255 4 1 3 3717 4193 3406 
0 4256 5 1 1 4194 
0 4257 4 1 3 3719 4195 3779 
0 4258 4 1 3 3720 4196 3780 
0 4283 7 1 2 4168 4036 
0 4284 7 2 2 4175 4037 
2 4285 1 4284  
2 4286 1 4284  
0 4287 3 3 2 3816 4238 
2 4288 1 4287  
2 4289 1 4287  
2 4290 1 4287  
0 4291 5 1 1 4187 
0 4295 5 1 1 4169 
0 4296 0 2 1 4170 
2 4297 1 4296  
2 4298 1 4296  
0 4299 5 1 1 4183 
0 4303 7 1 2 4252 2231 
0 4304 7 1 2 4256 2235 
0 4305 0 4 1 4198 
2 4306 1 4305  
2 4307 1 4305  
2 4308 1 4305  
2 4309 1 4305  
0 4310 3 3 2 3994 4283 
2 4311 1 4310  
2 4312 1 4310  
2 4313 1 4310  
0 4316 7 1 3 4176 4214 4204 
0 4317 7 1 2 4177 4210 
0 4318 7 1 3 4224 4131 4219 
0 4319 7 2 2 4225 4132 
2 4320 1 4319  
2 4321 1 4319  
0 4322 7 1 2 4171 4211 
0 4325 6 1 2 4205 3914 
0 4326 6 1 3 4206 4215 4172 
0 4327 6 1 2 4220 3817 
0 4328 6 1 3 4221 4133 3919 
0 4329 6 1 2 4248 4013 
0 4330 5 1 1 4249 
0 4331 7 2 3 334 4097 4295 
2 4332 1 4331  
2 4333 1 4331  
0 4335 7 2 2 4251 2730 
2 4336 1 4335  
2 4337 1 4335  
0 4338 7 2 2 4253 2734 
2 4339 1 4338  
2 4340 1 4338  
0 4341 7 2 2 4254 2736 
2 4342 1 4341  
2 4343 1 4341  
0 4344 7 2 2 4255 2738 
2 4345 1 4344  
2 4346 1 4344  
0 4347 7 2 2 4257 2742 
2 4348 1 4347  
2 4349 1 4347  
0 4350 7 2 2 4258 2744 
2 4351 1 4350  
2 4352 1 4350  
0 4353 0 2 1 4199 
2 4354 1 4353  
2 4355 1 4353  
0 4356 0 2 1 4207 
2 4357 1 4356  
2 4358 1 4356  
0 4359 0 2 1 4212 
2 4360 1 4359  
2 4361 1 4359  
0 4362 0 2 1 4222 
2 4363 1 4362  
2 4364 1 4362  
0 4365 0 2 1 4243 
2 4366 1 4365  
2 4367 1 4365  
0 4368 0 2 1 4244 
2 4369 1 4368  
2 4370 1 4368  
0 4371 7 2 2 4226 4227 
2 4372 1 4371  
2 4373 1 4371  
0 4376 4 1 3 3714 4303 2899 
0 4377 4 1 3 3718 4304 3642 
0 4387 7 2 2 335 4317 
2 4388 1 4387  
2 4389 1 4387  
0 4390 7 2 2 336 4318 
2 4391 1 4390  
2 4392 1 4390  
0 4393 6 1 2 3923 4330 
0 4398 0 2 1 4288 
2 4399 1 4398  
2 4400 1 4398  
0 4413 0 2 1 4285 
2 4414 1 4413  
2 4415 1 4413  
0 4416 6 2 3 3920 4325 4326 
2 4417 1 4416  
2 4418 1 4416  
0 4421 3 2 2 3814 4322 
2 4422 1 4421  
2 4423 1 4421  
0 4427 6 2 3 3948 4327 4328 
2 4428 1 4427  
2 4429 1 4427  
0 4430 0 2 1 4289 
2 4431 1 4430  
2 4432 1 4430  
0 4435 7 2 2 337 4316 
2 4436 1 4435  
2 4437 1 4435  
0 4442 3 1 2 4332 4297 
0 4443 7 2 4 4178 4306 4208 4216 
2 4444 1 4443  
2 4445 1 4443  
0 4446 6 1 2 4307 3811 
0 4447 6 1 3 4308 4201 3915 
0 4448 6 1 4 4309 4202 4217 4173 
0 4452 5 1 1 4357 
0 4458 6 2 2 4329 4393 
2 4459 1 4458  
2 4460 1 4458  
0 4461 5 1 1 4366 
0 4462 5 1 1 4369 
0 4463 6 1 2 4372 1460 
0 4464 5 1 1 4373 
0 4465 0 2 1 4311 
2 4466 1 4465  
2 4467 1 4465  
0 4468 4 2 2 4333 4298 
2 4469 1 4468  
2 4470 1 4468  
0 4472 7 2 2 4376 2732 
2 4473 1 4472  
2 4474 1 4472  
0 4475 7 2 2 4377 2740 
2 4476 1 4475  
2 4477 1 4475  
0 4479 0 2 1 4312 
2 4480 1 4479  
2 4481 1 4479  
0 4484 5 1 1 4354 
0 4486 5 1 1 4360 
0 4487 6 1 2 4361 4299 
0 4491 5 1 1 4363 
0 4493 7 2 2 338 4320 
2 4494 1 4493  
2 4495 1 4493  
0 4496 5 1 1 4399 
0 4497 7 1 2 4290 4400 
0 4498 7 2 2 4442 1769 
2 4499 1 4498  
2 4500 1 4498  
0 4503 6 2 4 3947 4446 4447 4448 
2 4504 1 4503  
2 4505 1 4503  
0 4506 5 1 1 4414 
0 4507 5 1 1 4436 
0 4508 5 1 1 4422 
0 4509 6 1 2 4423 4452 
0 4510 5 1 1 4428 
0 4511 6 1 2 4429 4241 
0 4515 6 1 2 967 4464 
0 4526 5 1 1 4417 
0 4527 6 1 2 4418 4484 
0 4528 6 1 2 4184 4486 
0 4529 5 1 1 4431 
0 4530 6 1 2 4432 4491 
0 4531 0 2 1 4388 
2 4532 1 4531  
2 4533 1 4531  
0 4534 0 2 1 4389 
2 4535 1 4534  
2 4536 1 4534  
0 4537 0 2 1 4391 
2 4538 1 4537  
2 4539 1 4537  
0 4540 0 2 1 4392 
2 4541 1 4540  
2 4542 1 4540  
0 4545 7 1 3 339 4321 4496 
0 4549 7 2 2 340 4444 
2 4550 1 4549  
2 4551 1 4549  
0 4552 6 1 2 4358 4508 
0 4555 6 1 2 4144 4510 
0 4558 5 1 1 4494 
0 4559 6 2 2 4463 4515 
2 4560 1 4559  
2 4561 1 4559  
0 4562 5 1 1 4466 
0 4563 7 1 2 4313 4467 
0 4564 0 3 1 4469 
2 4565 1 4564  
2 4566 1 4564  
2 4567 1 4564  
0 4568 5 1 1 4480 
0 4569 0 2 1 4445 
2 4570 1 4569  
2 4571 1 4569  
0 4572 6 1 2 4355 4526 
0 4573 6 1 2 4364 4529 
0 4576 6 2 2 4487 4528 
2 4577 1 4576  
2 4578 1 4576  
0 4581 0 2 1 4459 
2 4582 1 4581  
2 4583 1 4581  
0 4584 0 2 1 4460 
2 4585 1 4584  
2 4586 1 4584  
0 4587 3 1 3 2759 4499 2762 
0 4588 4 1 3 2760 4500 2763 
3 4589 3 0 2 4545 4497 
0 4593 6 2 2 4552 4509 
2 4594 1 4593  
2 4595 1 4593  
0 4596 5 1 1 4532 
0 4597 5 1 1 4535 
0 4599 6 2 2 4555 4511 
2 4600 1 4599  
2 4601 1 4599  
0 4602 5 1 1 4538 
0 4603 5 1 1 4541 
0 4608 7 1 3 341 4286 4562 
0 4613 0 2 1 4504 
2 4614 1 4613  
2 4615 1 4613  
0 4616 0 2 1 4505 
2 4617 1 4616  
2 4618 1 4616  
0 4619 6 2 2 4572 4527 
2 4620 1 4619  
2 4621 1 4619  
0 4623 6 2 2 4573 4530 
2 4624 1 4623  
2 4625 1 4623  
0 4628 5 1 1 4588 
0 4629 6 1 2 4570 4506 
0 4630 5 1 1 4571 
0 4635 5 1 1 4577 
0 4636 6 1 2 4578 4291 
0 4640 5 1 1 4582 
0 4641 6 1 2 4583 4461 
0 4642 5 1 1 4585 
0 4643 6 1 2 4586 4462 
0 4644 4 2 2 4608 4563 
2 4645 1 4644  
2 4646 1 4644  
0 4647 7 2 2 4560 2128 
2 4648 1 4647  
2 4649 1 4647  
0 4650 7 2 2 4561 2743 
2 4651 1 4650  
2 4652 1 4650  
0 4656 0 2 1 4550 
2 4657 1 4656  
2 4658 1 4656  
0 4659 0 2 1 4551 
2 4660 1 4659  
2 4661 1 4659  
0 4664 0 2 1 4565 
2 4665 1 4664  
2 4666 1 4664  
3 4667 7 0 2 4587 4628 
0 4668 6 1 2 4415 4630 
0 4669 5 1 1 4617 
0 4670 6 1 2 4618 4239 
0 4673 5 1 1 4620 
0 4674 6 1 2 4621 4507 
0 4675 6 1 2 4188 4635 
0 4676 5 1 1 4624 
0 4677 6 1 2 4625 4558 
0 4678 6 1 2 4367 4640 
0 4679 6 1 2 4370 4642 
0 4687 5 1 1 4614 
0 4688 6 1 2 4615 4568 
0 4691 0 2 1 4594 
2 4692 1 4691  
2 4693 1 4691  
0 4694 0 2 1 4595 
2 4695 1 4694  
2 4696 1 4694  
0 4697 0 2 1 4600 
2 4698 1 4697  
2 4699 1 4697  
0 4700 0 2 1 4601 
2 4701 1 4700  
2 4702 1 4700  
0 4704 6 1 2 4629 4668 
0 4705 6 1 2 4141 4669 
0 4706 5 1 1 4657 
0 4707 5 1 1 4660 
0 4708 6 1 2 4437 4673 
0 4711 6 2 2 4675 4636 
2 4712 1 4711  
2 4713 1 4711  
0 4716 6 1 2 4495 4676 
0 4717 6 3 2 4678 4641 
2 4718 1 4717  
2 4719 1 4717  
2 4720 1 4717  
0 4721 6 1 2 4679 4643 
0 4722 0 3 1 4645 
2 4723 1 4722  
2 4724 1 4722  
2 4725 1 4722  
0 4726 5 1 1 4665 
0 4727 3 2 3 4648 4651 4351 
2 4728 1 4727  
2 4729 1 4727  
0 4730 4 2 3 4649 4652 4352 
2 4731 1 4730  
2 4732 1 4730  
0 4733 6 1 2 4481 4687 
0 4740 6 2 2 4705 4670 
2 4741 1 4740  
2 4742 1 4740  
0 4743 6 3 2 4708 4674 
2 4744 1 4743  
2 4745 1 4743  
2 4746 1 4743  
0 4747 5 1 1 4692 
0 4748 6 1 2 4693 4596 
0 4749 5 1 1 4695 
0 4750 6 1 2 4696 4597 
0 4753 5 1 1 4698 
0 4754 6 1 2 4699 4602 
0 4755 5 1 1 4701 
0 4756 6 1 2 4702 4603 
0 4757 6 3 2 4716 4677 
2 4758 1 4757  
2 4759 1 4757  
2 4760 1 4757  
0 4769 6 2 2 4733 4688 
2 4770 1 4769  
2 4771 1 4769  
0 4772 7 2 2 342 4704 
2 4773 1 4772  
2 4774 1 4772  
0 4775 5 2 1 4721 
2 4776 1 4775  
2 4777 1 4775  
0 4778 5 1 1 4731 
0 4786 6 1 2 4533 4747 
0 4787 6 1 2 4536 4749 
0 4788 6 1 2 4539 4753 
0 4789 6 1 2 4542 4755 
0 4794 7 2 2 4712 2124 
2 4795 1 4794  
2 4796 1 4794  
0 4797 7 2 2 4713 2735 
2 4798 1 4797  
2 4799 1 4797  
0 4800 7 2 2 4718 2127 
2 4801 1 4800  
2 4802 1 4800  
0 4805 0 2 1 4723 
2 4806 1 4805  
2 4807 1 4805  
0 4808 7 2 2 4719 4470 
2 4809 1 4808  
2 4810 1 4808  
0 4812 0 2 1 4728 
2 4813 1 4812  
2 4814 1 4812  
3 4815 7 0 2 4729 4778 
0 4816 5 1 1 4770 
0 4817 5 1 1 4773 
0 4818 6 3 2 4786 4748 
2 4819 1 4818  
2 4820 1 4818  
2 4821 1 4818  
0 4822 6 1 2 4787 4750 
0 4823 6 2 2 4788 4754 
2 4824 1 4823  
2 4825 1 4823  
0 4826 6 1 2 4789 4756 
0 4829 6 1 2 4776 4726 
0 4830 5 1 1 4777 
0 4831 7 2 2 4744 2122 
2 4832 1 4831  
2 4833 1 4831  
0 4838 7 2 2 4758 2126 
2 4839 1 4838  
2 4840 1 4838  
0 4844 0 2 1 4741 
2 4845 1 4844  
2 4846 1 4844  
0 4847 0 2 1 4742 
2 4848 1 4847  
2 4849 1 4847  
0 4850 0 2 1 4745 
2 4851 1 4850  
2 4852 1 4850  
0 4854 0 2 1 4759 
2 4855 1 4854  
2 4856 1 4854  
0 4859 6 1 2 4774 4816 
0 4860 6 1 2 4771 4817 
0 4868 5 1 1 4826 
0 4870 5 1 1 4806 
0 4872 5 1 1 4809 
0 4873 6 1 2 4666 4830 
0 4876 3 3 3 4795 4798 4342 
2 4877 1 4876  
2 4878 1 4876  
2 4879 1 4876  
0 4880 4 2 3 4796 4799 4343 
2 4881 1 4880  
2 4882 1 4880  
0 4885 5 1 1 4813 
0 4889 5 2 1 4822 
2 4890 1 4889  
2 4891 1 4889  
0 4895 6 1 2 4859 4860 
0 4896 5 1 1 4845 
0 4897 6 1 2 4846 4706 
0 4898 5 1 1 4848 
0 4899 6 1 2 4849 4707 
0 4900 4 1 2 4868 4566 
0 4901 7 1 4 4720 4760 4824 4567 
0 4902 5 1 1 4851 
0 4904 5 1 1 4855 
0 4905 6 1 2 4856 4872 
0 4906 6 1 2 4873 4829 
0 4907 7 2 2 4819 2123 
2 4908 1 4907  
2 4909 1 4907  
0 4913 7 2 2 4825 2125 
2 4914 1 4913  
2 4915 1 4913  
0 4916 7 2 2 4820 4646 
2 4917 1 4916  
2 4918 1 4916  
0 4920 5 1 1 4881 
0 4921 7 2 2 4895 2184 
2 4922 1 4921  
2 4923 1 4921  
0 4924 6 1 2 4658 4896 
0 4925 6 1 2 4661 4898 
0 4926 3 1 2 4900 4901 
0 4928 6 1 2 4890 4870 
0 4929 5 1 1 4891 
0 4930 6 1 2 4810 4904 
0 4931 5 1 1 4906 
0 4937 0 2 1 4877 
2 4938 1 4937  
2 4939 1 4937  
0 4940 0 2 1 4878 
2 4941 1 4940  
2 4942 1 4940  
3 4944 7 0 2 4879 4920 
0 4946 6 2 2 4924 4897 
2 4947 1 4946  
2 4948 1 4946  
0 4949 6 1 2 4925 4899 
0 4950 6 1 2 4917 4902 
0 4951 5 1 1 4918 
0 4952 6 1 2 4807 4929 
0 4953 6 1 2 4930 4905 
0 4954 7 2 2 4926 2737 
2 4955 1 4954  
2 4956 1 4954  
0 4957 7 2 2 4931 2741 
2 4958 1 4957  
2 4959 1 4957  
0 4964 3 1 3 2765 2484 4922 
0 4965 4 1 3 2766 2485 4923 
0 4968 5 1 1 4949 
0 4969 6 1 2 4852 4951 
0 4970 6 1 2 4952 4928 
0 4973 7 2 2 4953 2739 
2 4974 1 4973  
2 4975 1 4973  
0 4978 5 1 1 4938 
0 4979 5 1 1 4941 
0 4980 5 1 1 4965 
0 4981 4 1 2 4968 4724 
0 4982 7 1 4 4821 4746 4947 4725 
0 4983 6 1 2 4950 4969 
0 4984 5 1 1 4970 
0 4985 7 2 2 4948 2121 
2 4986 1 4985  
2 4987 1 4985  
0 4988 3 2 3 4914 4955 4345 
2 4989 1 4988  
2 4990 1 4988  
0 4991 4 2 3 4915 4956 4346 
2 4992 1 4991  
2 4993 1 4991  
0 4996 3 2 3 4801 4958 4348 
2 4997 1 4996  
2 4998 1 4996  
0 4999 4 2 3 4802 4959 4349 
2 5000 1 4999  
2 5001 1 4999  
3 5002 7 0 2 4964 4980 
0 5007 3 1 2 4981 4982 
0 5010 7 2 2 4983 2731 
2 5011 1 5010  
2 5012 1 5010  
0 5013 7 2 2 4984 2733 
2 5014 1 5013  
2 5015 1 5013  
0 5018 3 2 3 4839 4974 4476 
2 5019 1 5018  
2 5020 1 5018  
0 5021 4 2 3 4840 4975 4477 
2 5022 1 5021  
2 5023 1 5021  
0 5026 5 1 1 4992 
0 5029 5 1 1 5000 
0 5030 7 2 2 5007 2729 
2 5031 1 5030  
2 5032 1 5030  
0 5039 0 2 1 4997 
2 5040 1 5039  
2 5041 1 5039  
0 5042 0 2 1 4989 
2 5043 1 5042  
2 5044 1 5042  
3 5045 7 0 2 4990 5026 
0 5046 5 1 1 5022 
3 5047 7 0 2 4998 5029 
0 5050 3 4 3 4832 5011 4473 
2 5051 1 5050  
2 5052 1 5050  
2 5053 1 5050  
2 5054 1 5050  
0 5055 4 2 3 4833 5012 4474 
2 5056 1 5055  
2 5057 1 5055  
0 5058 3 2 3 4908 5014 4339 
2 5059 1 5058  
2 5060 1 5058  
0 5061 4 2 3 4909 5015 4340 
2 5062 1 5061  
2 5063 1 5061  
0 5066 7 2 4 4732 5001 5023 4993 
2 5067 1 5066  
2 5068 1 5066  
0 5070 0 2 1 5019 
2 5071 1 5070  
2 5072 1 5070  
3 5078 7 0 2 5020 5046 
0 5080 3 4 3 4986 5031 4336 
2 5081 1 5080  
2 5082 1 5080  
2 5083 1 5080  
2 5084 1 5080  
0 5085 4 2 3 4987 5032 4337 
2 5086 1 5085  
2 5087 1 5085  
0 5094 6 1 2 5040 4885 
0 5095 5 1 1 5041 
0 5097 5 1 1 5043 
3 5102 7 0 2 5051 5052 
0 5103 5 1 1 5062 
0 5108 6 1 2 4814 5095 
0 5109 5 1 1 5071 
0 5110 6 1 2 5072 5097 
0 5111 0 2 1 5059 
2 5112 1 5111  
2 5113 1 5111  
0 5114 7 2 2 5053 1462 
2 5115 1 5114  
2 5116 1 5114  
0 5117 0 2 1 5054 
2 5118 1 5117  
2 5119 1 5117  
3 5120 7 0 2 5081 5082 
3 5121 7 0 2 5060 5103 
0 5122 6 2 2 5094 5108 
2 5123 1 5122  
2 5124 1 5122  
0 5125 6 1 2 5044 5109 
0 5128 7 2 2 1463 5083 
2 5129 1 5128  
2 5130 1 5128  
0 5133 7 2 4 4882 5063 5056 5086 
2 5134 1 5133  
2 5135 1 5133  
0 5136 7 1 3 5057 5087 1466 
0 5139 0 2 1 5084 
2 5140 1 5139  
2 5141 1 5139  
0 5145 6 2 2 5125 5110 
2 5146 1 5145  
2 5147 1 5145  
0 5151 0 2 1 5112 
2 5152 1 5151  
2 5153 1 5151  
0 5154 0 2 1 5113 
2 5155 1 5154  
2 5156 1 5154  
0 5159 5 1 1 5118 
0 5160 0 2 1 5115 
2 5161 1 5160  
2 5162 1 5160  
0 5163 0 2 1 5116 
2 5164 1 5163  
2 5165 1 5163  
0 5166 7 1 2 5067 5134 
0 5173 7 1 2 5068 5135 
0 5174 0 2 1 5123 
2 5175 1 5174  
2 5176 1 5174  
0 5177 0 2 1 5124 
2 5178 1 5177  
2 5179 1 5177  
0 5182 5 1 1 5140 
0 5183 6 1 2 5141 5159 
0 5184 0 2 1 5129 
2 5185 1 5184  
2 5186 1 5184  
0 5188 0 2 1 5130 
2 5189 1 5188  
2 5190 1 5188  
3 5192 5 0 1 5166 
0 5193 4 1 2 5136 5173 
0 5196 6 1 2 5152 4978 
0 5197 5 1 1 5153 
0 5198 6 1 2 5155 4979 
0 5199 5 1 1 5156 
0 5201 5 1 1 5161 
0 5203 5 1 1 5164 
0 5205 0 2 1 5146 
2 5206 1 5205  
2 5207 1 5205  
0 5209 0 2 1 5147 
2 5210 1 5209  
2 5211 1 5209  
0 5212 6 1 2 5119 5182 
0 5215 7 1 2 221 5193 
0 5217 5 1 1 5175 
0 5219 5 1 1 5178 
0 5220 6 1 2 4939 5197 
0 5221 6 1 2 4942 5199 
0 5222 5 1 1 5185 
0 5223 6 1 2 5186 5201 
0 5224 6 1 2 5189 5203 
0 5225 5 1 1 5190 
0 5228 6 2 2 5183 5212 
2 5229 1 5228  
2 5230 1 5228  
3 5231 5 0 1 5215 
0 5232 6 1 2 5206 5217 
0 5233 5 1 1 5207 
0 5234 6 1 2 5210 5219 
0 5235 5 1 1 5211 
0 5236 6 3 2 5196 5220 
2 5237 1 5236  
2 5238 1 5236  
2 5239 1 5236  
0 5240 6 1 2 5198 5221 
0 5242 6 1 2 5162 5222 
0 5243 6 1 2 5165 5225 
0 5245 6 1 2 5176 5233 
0 5246 6 1 2 5179 5235 
0 5250 5 2 1 5240 
2 5251 1 5250  
2 5252 1 5250  
0 5253 5 1 1 5229 
0 5254 6 2 2 5242 5223 
2 5255 1 5254  
2 5256 1 5254  
0 5257 6 1 2 5243 5224 
0 5258 6 2 2 5232 5245 
2 5259 1 5258  
2 5260 1 5258  
0 5261 6 1 2 5234 5246 
0 5266 5 2 1 5257 
2 5267 1 5266  
2 5268 1 5266  
0 5269 0 2 1 5237 
2 5270 1 5269  
2 5271 1 5269  
0 5277 7 1 3 5238 5255 2308 
0 5278 7 1 3 5251 5256 2311 
0 5279 5 2 1 5261 
2 5280 1 5279  
2 5281 1 5279  
0 5283 5 1 1 5270 
0 5284 6 1 2 5271 5253 
0 5285 7 1 3 5239 5267 2312 
0 5286 7 1 3 5252 5268 2309 
0 5289 0 2 1 5259 
2 5290 1 5289  
2 5291 1 5289  
0 5292 0 2 1 5260 
2 5293 1 5292  
2 5294 1 5292  
0 5295 6 1 2 5230 5283 
0 5298 3 2 4 5277 5285 5278 5286 
2 5299 1 5298  
2 5300 1 5298  
0 5303 0 2 1 5280 
2 5304 1 5303  
2 5305 1 5303  
0 5306 0 2 1 5281 
2 5307 1 5306  
2 5308 1 5306  
0 5309 6 2 2 5295 5284 
2 5310 1 5309  
2 5311 1 5309  
0 5312 5 1 1 5293 
0 5313 5 1 1 5290 
0 5322 5 1 1 5307 
0 5323 5 1 1 5304 
0 5324 0 2 1 5299 
2 5325 1 5324  
2 5326 1 5324  
0 5327 0 2 1 5300 
2 5328 1 5327  
2 5329 1 5327  
0 5332 0 2 1 5310 
2 5333 1 5332  
2 5334 1 5332  
0 5335 0 2 1 5311 
2 5336 1 5335  
2 5337 1 5335  
0 5340 6 1 2 5325 5323 
0 5341 6 1 2 5328 5322 
0 5344 5 1 1 5329 
0 5345 5 1 1 5326 
0 5348 6 1 2 5333 5313 
0 5349 6 1 2 5336 5312 
0 5350 6 1 2 5305 5345 
0 5351 6 1 2 5308 5344 
0 5352 5 1 1 5337 
0 5353 5 1 1 5334 
0 5354 6 1 2 5291 5353 
0 5355 6 1 2 5294 5352 
0 5356 6 1 2 5350 5340 
0 5357 6 1 2 5351 5341 
0 5358 6 1 2 5348 5354 
0 5359 6 1 2 5349 5355 
3 5360 7 0 2 5356 5357 
3 5361 6 0 2 5358 5359 
