1 1 0 2 0 
2 2 1 1  
2 3 1 1  
1 4 0 2 0 
2 5 1 4  
2 6 1 4  
0 2052 6 2 2 2036 2014 
2 2053 1 2052  
2 2054 1 2052  
1 7 0 2 0 
2 8 1 7  
2 9 1 7  
0 2055 6 2 2 2037 2016 
2 2056 1 2055  
2 2057 1 2055  
1 10 0 2 0 
2 11 1 10  
2 12 1 10  
0 2060 5 1 1 2038 
1 13 0 2 0 
2 14 1 13  
2 15 1 13  
0 2061 6 1 2 2039 2022 
0 2062 6 2 2 2040 294 
2 2063 1 2062  
2 2064 1 2062  
1 16 0 2 0 
2 17 1 16  
2 18 1 16  
1 19 0 2 0 
2 20 1 19  
2 21 1 19  
0 2067 5 1 1 2041 
0 2068 5 2 1 2028 
2 2069 1 2068  
2 2070 1 2068  
1 22 0 2 0 
2 23 1 22  
2 24 1 22  
0 2071 0 2 1 2029 
2 2072 1 2071  
2 2073 1 2071  
1 25 0 2 0 
2 26 1 25  
2 27 1 25  
1 28 0 2 0 
2 29 1 28  
2 30 1 28  
0 2076 5 1 1 2053 
0 2077 5 1 1 2056 
1 31 0 2 0 
2 32 1 31  
2 33 1 31  
0 2078 6 2 2 2060 295 
2 2079 1 2078  
2 2080 1 2078  
0 2081 6 2 2 2061 296 
2 2082 1 2081  
2 2083 1 2081  
1 34 0 2 0 
2 35 1 34  
2 36 1 34  
1 37 0 2 0 
2 38 1 37  
2 39 1 37  
0 2086 5 2 1 2043 
2 2087 1 2086  
2 2088 1 2086  
1 40 0 2 0 
2 41 1 40  
2 42 1 40  
0 2089 0 2 1 2044 
2 2090 1 2089  
2 2091 1 2089  
1 43 0 2 0 
2 44 1 43  
2 45 1 43  
1 46 0 2 0 
2 47 1 46  
2 48 1 46  
1 49 0 3 0 
2 50 1 49  
2 51 1 49  
2 52 1 49  
1 53 0 2 0 
2 54 1 53  
2 55 1 53  
1 56 0 3 0 
2 57 1 56  
2 58 1 56  
2 59 1 56  
0 2104 7 14 2 2031 2069 
2 2105 1 2104  
2 2106 1 2104  
2 2107 1 2104  
2 2108 1 2104  
2 2109 1 2104  
2 2110 1 2104  
2 2111 1 2104  
2 2112 1 2104  
2 2113 1 2104  
2 2114 1 2104  
2 2115 1 2104  
2 2116 1 2104  
2 2117 1 2104  
2 2118 1 2104  
1 60 0 2 0 
2 61 1 60  
2 62 1 60  
1 63 0 2 0 
2 64 1 63  
2 65 1 63  
1 66 0 2 0 
2 67 1 66  
2 68 1 66  
1 69 0 2 0 
2 70 1 69  
2 71 1 69  
0 2119 7 9 2 2034 2070 
2 2120 1 2119  
2 2121 1 2119  
2 2122 1 2119  
2 2123 1 2119  
2 2124 1 2119  
2 2125 1 2119  
2 2126 1 2119  
2 2127 1 2119  
2 2128 1 2119  
1 72 0 3 0 
2 73 1 72  
2 74 1 72  
2 75 1 72  
1 76 0 2 0 
2 77 1 76  
2 78 1 76  
1 79 0 2 0 
2 80 1 79  
2 81 1 79  
0 2129 7 13 2 2032 2072 
2 2130 1 2129  
2 2131 1 2129  
2 2132 1 2129  
2 2133 1 2129  
2 2134 1 2129  
2 2135 1 2129  
2 2136 1 2129  
2 2137 1 2129  
2 2138 1 2129  
2 2139 1 2129  
2 2140 1 2129  
2 2141 1 2129  
2 2142 1 2129  
1 82 0 2 0 
2 83 1 82  
2 84 1 82  
1 85 0 2 0 
2 86 1 85  
2 87 1 85  
1 88 0 2 0 
2 89 1 88  
2 90 1 88  
1 91 0 2 0 
2 92 1 91  
2 93 1 91  
1 94 0 4 0 
2 95 1 94  
2 96 1 94  
2 97 1 94  
2 98 1 94  
0 2143 7 4 2 2035 2073 
2 2144 1 2143  
2 2145 1 2143  
2 2146 1 2143  
2 2147 1 2143  
1 99 0 4 0 
2 100 1 99  
2 101 1 99  
2 102 1 99  
2 103 1 99  
0 2148 0 2 1 2063 
2 2149 1 2148  
2 2150 1 2148  
0 2151 0 2 1 2064 
2 2152 1 2151  
2 2153 1 2151  
1 104 0 7 0 
2 105 1 104  
2 106 1 104  
2 107 1 104  
2 108 1 104  
2 109 1 104  
2 110 1 104  
2 111 1 104  
0 2196 0 2 1 2079 
2 2197 1 2196  
2 2198 1 2196  
0 2199 0 2 1 2080 
2 2200 1 2199  
2 2201 1 2199  
0 2202 0 2 1 2082 
2 2203 1 2202  
2 2204 1 2202  
0 2205 0 2 1 2083 
2 2206 1 2205  
2 2207 1 2205  
0 2214 6 1 2 2152 915 
0 2215 5 1 1 2153 
0 2216 6 1 2 2149 916 
0 2217 5 1 1 2150 
0 2222 6 1 2 2200 1348 
0 2223 5 1 1 2201 
0 2224 6 1 2 2197 1349 
0 2225 5 1 1 2198 
0 2226 6 1 2 2206 913 
0 2227 5 1 1 2207 
0 2228 6 1 2 2203 914 
0 2229 5 1 1 2204 
0 2230 6 1 2 669 2215 
0 2231 6 1 2 666 2217 
0 2232 6 1 2 1257 2223 
0 2233 6 1 2 1254 2225 
0 2234 6 1 2 663 2227 
0 2235 6 1 2 660 2229 
0 2236 6 1 2 2214 2230 
0 2237 6 2 2 2216 2231 
2 2238 1 2237  
2 2239 1 2237  
0 190 5 3 1 2 
2 191 1 190  
2 192 1 190  
2 193 1 190  
0 2240 6 1 2 2222 2232 
0 2241 6 2 2 2224 2233 
2 2242 1 2241  
2 2243 1 2241  
0 194 5 2 1 5 
2 195 1 194  
2 196 1 194  
0 2244 6 1 2 2226 2234 
0 197 5 3 1 8 
2 198 1 197  
2 199 1 197  
2 200 1 197  
0 2245 6 2 2 2228 2235 
2 2246 1 2245  
2 2247 1 2245  
0 201 5 4 1 11 
2 202 1 201  
2 203 1 201  
2 204 1 201  
2 205 1 201  
0 2250 5 1 1 2236 
0 2253 5 1 1 2240 
0 206 5 2 1 14 
2 207 1 206  
2 208 1 206  
0 2256 5 1 1 2244 
0 209 5 2 1 17 
2 210 1 209  
2 211 1 209  
0 2257 5 2 1 2238 
2 2258 1 2257  
2 2259 1 2257  
0 212 5 3 1 20 
2 213 1 212  
2 214 1 212  
2 215 1 212  
0 2260 0 2 1 2239 
2 2261 1 2260  
2 2262 1 2260  
0 2263 5 2 1 2242 
2 2264 1 2263  
2 2265 1 2263  
0 216 5 3 1 23 
2 217 1 216  
2 218 1 216  
2 219 1 216  
0 2266 7 2 2 1165 2243 
2 2267 1 2266  
2 2268 1 2266  
0 220 5 4 1 26 
2 221 1 220  
2 222 1 220  
2 223 1 220  
2 224 1 220  
0 2269 5 2 1 2246 
2 2270 1 2269  
2 2271 1 2269  
0 2272 7 2 2 1169 2247 
2 2273 1 2272  
2 2274 1 2272  
0 225 5 3 1 29 
2 226 1 225  
2 227 1 225  
2 228 1 225  
0 229 5 2 1 32 
2 230 1 229  
2 231 1 229  
0 2279 6 2 8 2067 2012 2047 2250 902 2256 2253 906 
2 2280 1 2279  
2 2281 1 2279  
0 232 5 2 1 35 
2 233 1 232  
2 234 1 232  
0 235 5 3 1 38 
2 236 1 235  
2 237 1 235  
2 238 1 235  
0 2286 0 10 1 2267 
2 2287 1 2286  
2 2288 1 2286  
2 2289 1 2286  
2 2290 1 2286  
2 2291 1 2286  
2 2292 1 2286  
2 2293 1 2286  
2 2294 1 2286  
2 2295 1 2286  
2 2296 1 2286  
0 239 5 3 1 41 
2 240 1 239  
2 241 1 239  
2 242 1 239  
0 243 5 3 1 44 
2 244 1 243  
2 245 1 243  
2 246 1 243  
0 247 5 3 1 47 
2 248 1 247  
2 249 1 247  
2 250 1 247  
0 2297 0 15 1 2268 
2 2298 1 2297  
2 2299 1 2297  
2 2300 1 2297  
2 2301 1 2297  
2 2302 1 2297  
2 2303 1 2297  
2 2304 1 2297  
2 2305 1 2297  
2 2306 1 2297  
2 2307 1 2297  
2 2308 1 2297  
2 2309 1 2297  
2 2310 1 2297  
2 2311 1 2297  
2 2312 1 2297  
0 251 6 1 2 64 89 
0 252 6 1 2 67 92 
0 253 5 2 1 73 
2 254 1 253  
2 255 1 253  
0 256 5 1 1 74 
0 257 0 2 1 70 
2 258 1 257  
2 259 1 257  
0 260 0 2 1 71 
2 261 1 260  
2 262 1 260  
0 263 5 2 1 77 
2 264 1 263  
2 265 1 263  
0 266 5 2 1 80 
2 267 1 266  
2 268 1 266  
0 2315 0 10 1 2273 
2 2316 1 2315  
2 2317 1 2315  
2 2318 1 2315  
2 2319 1 2315  
2 2320 1 2315  
2 2321 1 2315  
2 2322 1 2315  
2 2323 1 2315  
2 2324 1 2315  
2 2325 1 2315  
0 269 5 2 1 83 
2 270 1 269  
2 271 1 269  
0 272 5 2 1 86 
2 273 1 272  
2 274 1 272  
0 275 5 1 1 105 
0 276 5 1 1 106 
0 277 5 2 1 90 
2 278 1 277  
2 279 1 277  
0 2326 0 13 1 2274 
2 2327 1 2326  
2 2328 1 2326  
2 2329 1 2326  
2 2330 1 2326  
2 2331 1 2326  
2 2332 1 2326  
2 2333 1 2326  
2 2334 1 2326  
2 2335 1 2326  
2 2336 1 2326  
2 2337 1 2326  
2 2338 1 2326  
2 2339 1 2326  
0 280 5 2 1 93 
2 281 1 280  
2 282 1 280  
0 283 0 6 1 95 
2 284 1 283  
2 285 1 283  
2 286 1 283  
2 287 1 283  
2 288 1 283  
2 289 1 283  
0 290 5 6 1 96 
2 291 1 290  
2 292 1 290  
2 293 1 290  
2 294 1 290  
2 295 1 290  
2 296 1 290  
0 2340 7 12 2 2087 2258 
2 2341 1 2340  
2 2342 1 2340  
2 2343 1 2340  
2 2344 1 2340  
2 2345 1 2340  
2 2346 1 2340  
2 2347 1 2340  
2 2348 1 2340  
2 2349 1 2340  
2 2350 1 2340  
2 2351 1 2340  
2 2352 1 2340  
0 297 0 2 1 97 
2 298 1 297  
2 299 1 297  
0 300 5 2 1 98 
2 301 1 300  
2 302 1 300  
0 303 0 2 1 100 
2 304 1 303  
2 305 1 303  
0 2353 7 7 2 2090 2259 
2 2354 1 2353  
2 2355 1 2353  
2 2356 1 2353  
2 2357 1 2353  
2 2358 1 2353  
2 2359 1 2353  
2 2360 1 2353  
0 306 5 6 1 101 
2 307 1 306  
2 308 1 306  
2 309 1 306  
2 310 1 306  
2 311 1 306  
2 312 1 306  
0 313 5 2 1 102 
2 314 1 313  
2 315 1 313  
0 2361 7 13 2 2088 2261 
2 2362 1 2361  
2 2363 1 2361  
2 2364 1 2361  
2 2365 1 2361  
2 2366 1 2361  
2 2367 1 2361  
2 2368 1 2361  
2 2369 1 2361  
2 2370 1 2361  
2 2371 1 2361  
2 2372 1 2361  
2 2373 1 2361  
2 2374 1 2361  
0 316 0 2 1 107 
2 317 1 316  
2 318 1 316  
0 319 5 6 1 108 
2 320 1 319  
2 321 1 319  
2 322 1 319  
2 323 1 319  
2 324 1 319  
2 325 1 319  
0 326 0 4 1 109 
2 327 1 326  
2 328 1 326  
2 329 1 326  
2 330 1 326  
0 2375 7 8 2 2091 2262 
2 2376 1 2375  
2 2377 1 2375  
2 2378 1 2375  
2 2379 1 2375  
2 2380 1 2375  
2 2381 1 2375  
2 2382 1 2375  
2 2383 1 2375  
0 331 0 6 1 110 
2 332 1 331  
2 333 1 331  
2 334 1 331  
2 335 1 331  
2 336 1 331  
2 337 1 331  
0 2384 7 1 4 341 2280 314 315 
0 2385 7 1 2 1163 2264 
0 338 5 4 1 111 
2 339 1 338  
2 340 1 338  
2 341 1 338  
2 342 1 338  
0 2386 7 14 2 1166 2265 
2 2387 1 2386  
2 2388 1 2386  
2 2389 1 2386  
2 2390 1 2386  
2 2391 1 2386  
2 2392 1 2386  
2 2393 1 2386  
2 2394 1 2386  
2 2395 1 2386  
2 2396 1 2386  
2 2397 1 2386  
2 2398 1 2386  
2 2399 1 2386  
2 2400 1 2386  
0 343 0 2 1 3 
2 344 1 343  
2 345 1 343  
0 346 0 2 1 6 
2 347 1 346  
2 348 1 346  
0 349 0 2 1 9 
2 350 1 349  
2 351 1 349  
0 352 0 2 1 12 
2 353 1 352  
2 354 1 352  
0 355 0 2 1 15 
2 356 1 355  
2 357 1 355  
0 358 0 2 1 18 
2 359 1 358  
2 360 1 358  
0 361 0 2 1 21 
2 362 1 361  
2 363 1 361  
0 364 0 2 1 24 
2 365 1 364  
2 366 1 364  
0 367 0 2 1 27 
2 368 1 367  
2 369 1 367  
0 370 0 2 1 30 
2 371 1 370  
2 372 1 370  
0 373 0 2 1 33 
2 374 1 373  
2 375 1 373  
0 376 0 2 1 36 
2 377 1 376  
2 378 1 376  
0 2426 7 1 2 1167 2270 
0 379 0 2 1 39 
2 380 1 379  
2 381 1 379  
0 2427 7 16 2 1170 2271 
2 2428 1 2427  
2 2429 1 2427  
2 2430 1 2427  
2 2431 1 2427  
2 2432 1 2427  
2 2433 1 2427  
2 2434 1 2427  
2 2435 1 2427  
2 2436 1 2427  
2 2437 1 2427  
2 2438 1 2427  
2 2439 1 2427  
2 2440 1 2427  
2 2441 1 2427  
2 2442 1 2427  
2 2443 1 2427  
0 382 0 2 1 42 
2 383 1 382  
2 384 1 382  
0 385 0 2 1 45 
2 386 1 385  
2 387 1 385  
0 388 0 2 1 48 
2 389 1 388  
2 390 1 388  
0 2537 6 2 5 2287 2316 2362 2105 1172 
2 2538 1 2537  
2 2539 1 2537  
0 2540 6 2 5 2288 2317 2341 2130 1173 
2 2541 1 2540  
2 2542 1 2540  
0 2543 6 2 5 2289 2318 2342 2120 1174 
2 2544 1 2543  
2 2545 1 2543  
0 2546 6 2 5 2290 2319 2354 2106 1175 
2 2547 1 2546  
2 2548 1 2546  
0 2549 6 2 5 2298 2320 2376 2121 1189 
2 2550 1 2549  
2 2551 1 2549  
0 2552 6 2 5 2299 2327 2363 2144 1190 
2 2553 1 2552  
2 2554 1 2552  
0 2555 6 2 5 2300 2328 2377 2131 1191 
2 2556 1 2555  
2 2557 1 2555  
0 2558 7 2 5 2291 2321 2364 2107 1176 
2 2559 1 2558  
2 2560 1 2558  
0 2561 7 2 5 2292 2322 2343 2132 1177 
2 2562 1 2561  
2 2563 1 2561  
0 2564 7 2 5 2293 2323 2344 2122 1178 
2 2565 1 2564  
2 2566 1 2564  
0 2567 7 2 5 2294 2324 2355 2108 1179 
2 2568 1 2567  
2 2569 1 2567  
0 2570 7 2 5 2301 2325 2378 2123 1192 
2 2571 1 2570  
2 2572 1 2570  
0 2573 7 2 5 2302 2329 2365 2145 1193 
2 2574 1 2573  
2 2575 1 2573  
0 2576 7 2 5 2303 2330 2379 2133 1194 
2 2577 1 2576  
2 2578 1 2576  
0 534 5 1 1 344 
0 535 5 1 1 347 
0 536 5 1 1 350 
0 537 5 1 1 353 
0 538 5 1 1 356 
0 539 5 1 1 359 
0 540 5 1 1 362 
0 541 5 1 1 365 
0 542 5 1 1 368 
0 543 5 1 1 371 
0 544 5 1 1 374 
0 545 5 1 1 377 
0 546 5 1 1 380 
0 547 5 1 1 383 
0 548 5 1 1 386 
0 549 5 1 1 389 
0 550 6 1 2 307 332 
0 551 6 1 2 308 333 
0 552 6 1 2 309 334 
0 553 6 1 2 310 335 
0 554 6 1 2 311 336 
0 555 6 1 2 312 337 
0 556 0 2 1 191 
2 557 1 556  
2 558 1 556  
0 2597 6 2 5 2304 2429 2367 2124 1181 
2 2598 1 2597  
2 2599 1 2597  
0 2600 6 2 5 2305 2430 2380 2109 1182 
2 2601 1 2600  
2 2602 1 2600  
0 559 0 2 1 195 
2 560 1 559  
2 561 1 559  
0 2603 6 2 5 2306 2431 2345 2146 1183 
2 2604 1 2603  
2 2605 1 2603  
0 2606 6 2 5 2307 2432 2356 2135 1195 
2 2607 1 2606  
2 2608 1 2606  
0 562 0 2 1 207 
2 563 1 562  
2 564 1 562  
0 2611 6 2 5 2387 2331 2368 2136 1196 
2 2612 1 2611  
2 2613 1 2611  
0 565 0 2 1 210 
2 566 1 565  
2 567 1 565  
0 2614 6 2 5 2388 2332 2369 2125 1197 
2 2615 1 2614  
2 2616 1 2614  
0 568 0 2 1 226 
2 569 1 568  
2 570 1 568  
0 2617 6 2 5 2389 2333 2381 2110 1198 
2 2618 1 2617  
2 2619 1 2617  
0 571 0 2 1 244 
2 572 1 571  
2 573 1 571  
0 2620 6 2 5 2390 2334 2357 2137 1199 
2 2621 1 2620  
2 2622 1 2620  
0 574 7 2 2 65 320 
2 575 1 574  
2 576 1 574  
0 577 0 2 1 221 
2 578 1 577  
2 579 1 577  
0 2627 6 1 5 2308 2433 2346 2111 927 
0 580 0 2 1 230 
2 581 1 580  
2 582 1 580  
0 2628 6 1 5 2391 2335 2347 2112 928 
0 2629 6 1 5 2392 2434 2370 2113 929 
0 583 0 2 1 233 
2 584 1 583  
2 585 1 583  
0 2630 6 1 5 2393 2435 2348 2138 930 
0 2631 6 1 5 2394 2436 2349 2126 931 
0 586 7 2 2 68 321 
2 587 1 586  
2 588 1 586  
0 2632 6 1 5 2395 2437 2358 2114 932 
0 2633 6 1 5 2396 2426 2350 2115 933 
0 589 0 2 1 240 
2 590 1 589  
2 591 1 589  
0 2634 6 1 5 2385 2438 2351 2116 934 
0 2639 7 2 5 2296 2439 2371 2139 1184 
2 2640 1 2639  
2 2641 1 2639  
0 592 7 2 3 50 254 322 
2 593 1 592  
2 594 1 592  
0 2642 7 2 5 2309 2440 2372 2127 1185 
2 2643 1 2642  
2 2644 1 2642  
0 595 0 2 1 248 
2 596 1 595  
2 597 1 595  
0 2645 7 2 5 2310 2441 2382 2117 1186 
2 2646 1 2645  
2 2647 1 2645  
0 598 0 2 1 241 
2 599 1 598  
2 600 1 598  
0 2648 7 2 5 2311 2442 2352 2147 1187 
2 2649 1 2648  
2 2650 1 2648  
0 601 6 1 2 327 278 
0 602 6 1 2 328 281 
0 603 6 4 2 261 75 
2 604 1 603  
2 605 1 603  
2 606 1 603  
2 607 1 603  
0 2651 7 2 5 2312 2443 2359 2140 1200 
2 2652 1 2651  
2 2653 1 2651  
0 2655 7 2 5 2397 2336 2373 2141 1201 
2 2656 1 2655  
2 2657 1 2655  
0 608 6 3 2 262 301 
2 609 1 608  
2 610 1 608  
2 611 1 608  
0 2658 7 2 5 2398 2337 2374 2128 1202 
2 2659 1 2658  
2 2660 1 2658  
0 612 6 3 2 256 302 
2 613 1 612  
2 614 1 612  
2 615 1 612  
0 2661 7 2 5 2399 2338 2383 2118 1203 
2 2662 1 2661  
2 2663 1 2661  
0 616 0 2 1 202 
2 617 1 616  
2 618 1 616  
0 2664 7 2 5 2400 2339 2360 2142 1204 
2 2665 1 2664  
2 2666 1 2664  
0 619 0 2 1 217 
2 620 1 619  
2 621 1 619  
0 2669 6 1 2 2559 534 
0 622 0 2 1 222 
2 623 1 622  
2 624 1 622  
0 2670 5 1 1 2560 
0 2671 6 1 2 2562 535 
0 625 0 2 1 242 
2 626 1 625  
2 627 1 625  
0 2672 5 1 1 2563 
0 2673 6 1 2 2565 536 
0 628 0 2 1 192 
2 629 1 628  
2 630 1 628  
0 2674 5 1 1 2566 
0 2675 6 1 2 2568 537 
0 631 0 2 1 193 
2 632 1 631  
2 633 1 631  
0 2676 5 1 1 2569 
0 634 0 2 1 196 
2 635 1 634  
2 636 1 634  
0 2682 6 1 2 2571 543 
0 2683 5 1 1 2572 
0 637 0 2 1 231 
2 638 1 637  
2 639 1 637  
0 640 0 2 1 198 
2 641 1 640  
2 642 1 640  
0 2688 6 1 2 2574 548 
0 2689 5 1 1 2575 
0 643 7 2 3 57 258 323 
2 644 1 643  
2 645 1 643  
0 2690 6 1 2 2577 549 
0 2691 5 1 1 2578 
0 646 0 2 1 234 
2 647 1 646  
2 648 1 646  
0 649 0 2 1 203 
2 650 1 649  
2 651 1 649  
0 652 0 2 1 236 
2 653 1 652  
2 654 1 652  
0 655 7 2 3 61 259 324 
2 656 1 655  
2 657 1 655  
0 658 0 2 1 264 
2 659 1 658  
2 660 1 658  
0 661 0 2 1 265 
2 662 1 661  
2 663 1 661  
0 2710 7 1 8 2627 2628 2629 2630 2631 2632 2633 2634 
0 664 0 2 1 267 
2 665 1 664  
2 666 1 664  
0 667 0 2 1 268 
2 668 1 667  
2 669 1 667  
0 670 0 2 1 270 
2 671 1 670  
2 672 1 670  
0 2720 6 1 2 345 2670 
0 673 0 2 1 271 
2 674 1 673  
2 675 1 673  
0 2721 6 1 2 348 2672 
0 2722 6 1 2 351 2674 
0 676 0 2 1 273 
2 677 1 676  
2 678 1 676  
0 2723 6 1 2 354 2676 
0 2724 6 1 2 2640 538 
0 679 0 2 1 274 
2 680 1 679  
2 681 1 679  
0 2725 5 1 1 2641 
0 2726 6 1 2 2643 539 
0 682 7 2 2 251 317 
2 683 1 682  
2 684 1 682  
0 2727 5 1 1 2644 
0 2728 6 1 2 2646 540 
0 685 7 2 2 252 318 
2 686 1 685  
2 687 1 685  
0 2729 5 1 1 2647 
0 2730 6 1 2 2649 541 
0 688 0 2 1 199 
2 689 1 688  
2 690 1 688  
0 2731 5 1 1 2650 
0 2732 6 1 2 2652 542 
0 691 0 2 1 200 
2 692 1 691  
2 693 1 691  
0 2733 5 1 1 2653 
0 2734 6 1 2 372 2683 
0 694 0 2 1 213 
2 695 1 694  
2 696 1 694  
0 2735 6 1 2 2656 544 
0 2736 5 1 1 2657 
0 697 0 2 1 214 
2 698 1 697  
2 699 1 697  
0 2737 6 1 2 2659 545 
0 2738 5 1 1 2660 
0 700 0 2 1 249 
2 701 1 700  
2 702 1 700  
0 2740 5 1 1 2663 
0 2741 6 1 2 2665 547 
0 703 0 2 1 250 
2 704 1 703  
2 705 1 703  
0 2743 6 1 2 387 2689 
0 2744 6 1 2 390 2691 
0 706 0 2 1 237 
2 707 1 706  
2 708 1 706  
0 2746 6 1 8 2607 2550 2612 2615 2618 2621 2553 2556 
0 2747 7 2 8 2539 2542 2545 2548 2596 2599 2602 2605 
2 2748 1 2747  
2 2749 1 2747  
0 709 0 2 1 238 
2 710 1 709  
2 711 1 709  
0 2750 7 2 8 2608 2551 2613 2616 2619 2622 2554 2557 
2 2751 1 2750  
2 2752 1 2750  
3 2753 6 0 2 2669 2720 
0 712 0 2 1 204 
2 713 1 712  
2 714 1 712  
3 2754 6 0 2 2671 2721 
3 2755 6 0 2 2673 2722 
0 715 0 2 1 205 
2 716 1 715  
2 717 1 715  
3 2756 6 0 2 2675 2723 
0 2757 6 1 2 357 2725 
0 718 0 2 1 208 
2 719 1 718  
2 720 1 718  
0 2758 6 1 2 360 2727 
0 2759 6 1 2 363 2729 
0 721 0 2 1 218 
2 722 1 721  
2 723 1 721  
0 2761 6 1 2 369 2733 
3 2762 6 0 2 2682 2734 
0 724 7 2 3 54 255 325 
2 725 1 724  
2 726 1 724  
0 2764 6 1 2 378 2738 
0 2765 6 1 2 381 2740 
0 727 0 2 1 245 
2 728 1 727  
2 729 1 727  
3 2767 6 0 2 2688 2743 
3 2768 6 0 2 2690 2744 
2 730 0 2 1 223 
2 731 1 730  
2 732 1 730  
0 2773 7 2 2 2745 275 
0 2774 -1 1  
2 2775 1 2776  
2 2776 7 2 2 2746 276 
0 2777 -1 1  
0 2778 -1 1  
0 733 0 2 1 224 
2 734 1 733  
2 735 1 733  
3 2779 6 0 2 2724 2757 
3 2780 6 0 2 2726 2758 
0 736 0 2 1 211 
2 737 1 736  
2 738 1 736  
3 2781 6 0 2 2728 2759 
3 2782 6 0 2 2730 2760 
0 739 0 2 1 219 
2 740 1 739  
2 741 1 739  
3 2783 6 0 2 2732 2761 
3 2784 6 0 2 2735 2763 
0 742 0 2 1 227 
2 743 1 742  
2 744 1 742  
3 2785 6 0 2 2737 2764 
3 2786 6 0 2 2739 2765 
0 745 0 2 1 246 
2 746 1 745  
2 747 1 745  
3 2787 6 0 2 2741 2766 
2 2788 7 2789 3 2748 2751 2710 
2 748 0 2 1 215 
2 749 1 748  
2 750 1 748  
2 2789 6 6 2 2749 2752 
0 2790 -1 1  
0 2791 -1 1  
0 2792 -1 1  
0 2793 -1 1  
0 2794 -1 1  
0 2795 -1 1  
0 751 0 2 1 228 
2 752 1 751  
2 753 1 751  
0 2800 7 1 4 342 2281 103 2788 
0 2807 6 1 2 2774 2018 
0 2808 5 1 1 2775 
0 2809 6 1 2 2777 2019 
0 2810 5 1 1 2778 
3 2811 4 0 2 2384 2800 
0 2594 6 2 5 2295 2428 2366 2134 1180 
2 2595 1 2594  
2 2596 1 2594  
0 2812 7 2 3 897 284 2790 
2 2813 1 2812  
2 2814 1 2812  
0 2815 7 2 3 78 285 2791 
2 2816 1 2815  
2 2817 1 2815  
0 2818 7 2 3 84 286 2792 
2 2819 1 2818  
2 2820 1 2818  
0 2821 7 2 3 87 287 2793 
2 2822 1 2821  
2 2823 1 2821  
0 2824 7 2 3 898 288 2794 
2 2825 1 2824  
2 2826 1 2824  
0 2827 6 1 2 1967 2808 
0 2828 6 1 2 1970 2810 
0 2829 7 2 3 81 289 2795 
2 2830 1 2829  
2 2831 1 2829  
0 2843 6 2 2 2807 2827 
2 2844 1 2843  
2 2845 1 2843  
0 2846 6 2 2 2809 2828 
2 2847 1 2846  
2 2848 1 2846  
0 2850 6 1 2 2813 2076 
0 2851 6 1 2 2816 2077 
0 2852 6 1 2 2819 1915 
0 2853 6 1 2 2822 1857 
0 2854 6 1 2 2825 1938 
0 2857 5 1 1 2814 
0 2858 5 1 1 2817 
0 2859 5 1 1 2820 
0 2860 5 1 1 2823 
0 2861 5 1 1 2826 
0 2862 5 1 1 2830 
0 2863 6 1 2 2831 1985 
0 2866 6 1 2 2054 2857 
0 2867 6 1 2 2057 2858 
0 2868 6 1 2 1868 2859 
0 2869 6 1 2 1820 2860 
0 2870 6 1 2 1904 2861 
0 2871 6 1 2 2844 886 
0 2872 5 1 1 2845 
0 2873 6 1 2 2847 887 
0 2874 5 1 1 2848 
0 2875 6 1 2 1935 2862 
0 2876 6 1 2 2866 2850 
0 2877 6 1 2 2867 2851 
0 2878 6 1 2 2868 2852 
0 2879 6 1 2 2869 2853 
0 2880 6 1 2 2870 2854 
0 2881 6 1 2 684 2872 
0 2882 6 1 2 687 2874 
0 2883 6 2 2 2875 2863 
2 2884 1 2883  
2 2885 1 2883  
3 2886 7 0 2 2876 550 
3 2887 7 0 2 551 2877 
3 2888 7 0 2 553 2878 
3 2889 7 0 2 2879 554 
3 2890 7 0 2 555 2880 
3 2891 6 0 2 2871 2881 
3 2892 6 0 2 2873 2882 
0 2895 6 1 2 2884 1461 
0 2896 5 1 1 2885 
0 2897 6 1 2 1385 2896 
0 2898 6 1 2 2895 2897 
3 2899 7 0 2 2898 552 
0 886 5 1 1 683 
0 887 5 1 1 686 
0 888 5 1 1 617 
0 889 5 1 1 620 
0 890 5 1 1 623 
0 891 5 1 1 626 
0 892 5 1 1 632 
0 893 5 1 1 644 
0 894 5 1 1 650 
0 895 5 1 1 653 
0 896 5 1 1 656 
0 897 7 1 2 51 613 
0 898 7 1 2 58 609 
0 899 6 3 2 55 614 
2 900 1 899  
2 901 1 899  
2 902 1 899  
0 903 6 3 2 62 610 
2 904 1 903  
2 905 1 903  
2 906 1 903  
0 907 6 2 2 52 615 
2 908 1 907  
2 909 1 907  
0 910 6 2 2 59 611 
2 911 1 910  
2 912 1 910  
0 913 5 1 1 662 
0 914 5 1 1 659 
0 915 5 1 1 668 
0 916 5 1 1 665 
0 917 5 1 1 674 
0 918 5 1 1 671 
0 919 5 1 1 680 
0 920 5 1 1 677 
0 921 6 1 4 279 298 329 604 
0 922 6 1 4 282 299 330 605 
0 923 6 2 3 304 339 606 
2 924 1 923  
2 925 1 923  
0 926 7 8 3 305 340 607 
2 927 1 926  
2 928 1 926  
2 929 1 926  
2 930 1 926  
2 931 1 926  
2 932 1 926  
2 933 1 926  
2 934 1 926  
0 935 0 2 1 557 
2 936 1 935  
2 937 1 935  
0 938 5 1 1 689 
0 939 0 2 1 558 
2 940 1 939  
2 941 1 939  
0 942 5 1 1 692 
0 943 0 2 1 563 
2 944 1 943  
2 945 1 943  
0 946 5 1 1 695 
0 947 0 2 1 564 
2 948 1 947  
2 949 1 947  
0 950 5 1 1 698 
0 951 0 2 1 569 
2 952 1 951  
2 953 1 951  
0 954 5 1 1 701 
0 955 0 2 1 570 
2 956 1 955  
2 957 1 955  
0 958 5 1 1 704 
0 959 0 2 1 575 
2 960 1 959  
2 961 1 959  
0 962 0 2 1 576 
2 963 1 962  
2 964 1 962  
0 965 0 2 1 581 
2 966 1 965  
2 967 1 965  
0 968 5 1 1 707 
0 969 0 2 1 582 
2 970 1 969  
2 971 1 969  
0 972 5 1 1 710 
0 973 0 2 1 587 
2 974 1 973  
2 975 1 973  
0 976 5 1 1 713 
0 977 0 2 1 588 
2 978 1 977  
2 979 1 977  
0 980 5 1 1 716 
0 981 0 2 1 593 
2 982 1 981  
2 983 1 981  
0 984 5 1 1 629 
0 985 0 2 1 594 
2 986 1 985  
2 987 1 985  
0 988 5 1 1 719 
0 989 5 1 1 722 
0 990 5 1 1 635 
0 991 5 1 1 725 
0 992 5 1 1 728 
0 993 5 1 1 638 
0 994 0 2 1 596 
2 995 1 994  
2 996 1 994  
0 997 5 1 1 731 
0 998 0 2 1 597 
2 999 1 998  
2 1000 1 998  
0 1001 5 1 1 734 
0 1002 5 1 1 737 
0 1003 5 1 1 740 
0 1004 5 1 1 641 
0 1005 5 1 1 743 
0 1006 5 1 1 746 
0 1007 5 1 1 647 
0 1008 5 1 1 749 
0 1009 5 1 1 752 
0 1010 0 2 1 560 
2 1011 1 1010  
2 1012 1 1010  
0 1013 0 2 1 561 
2 1014 1 1013  
2 1015 1 1013  
0 1016 0 2 1 566 
2 1017 1 1016  
2 1018 1 1016  
0 1019 0 2 1 567 
2 1020 1 1019  
2 1021 1 1019  
0 1022 0 2 1 572 
2 1023 1 1022  
2 1024 1 1022  
0 1025 0 2 1 573 
2 1026 1 1025  
2 1027 1 1025  
0 1028 0 2 1 578 
2 1029 1 1028  
2 1030 1 1028  
0 1031 0 2 1 579 
2 1032 1 1031  
2 1033 1 1031  
0 1034 0 2 1 584 
2 1035 1 1034  
2 1036 1 1034  
0 1037 0 2 1 585 
2 1038 1 1037  
2 1039 1 1037  
0 1040 0 2 1 590 
2 1041 1 1040  
2 1042 1 1040  
0 1043 0 2 1 591 
2 1044 1 1043  
2 1045 1 1043  
0 1046 0 2 1 599 
2 1047 1 1046  
2 1048 1 1046  
0 1049 0 2 1 600 
2 1050 1 1049  
2 1051 1 1049  
0 1054 6 1 2 621 888 
0 1055 6 1 2 618 889 
0 1063 6 1 2 627 890 
0 1064 6 1 2 624 891 
0 1067 6 1 2 657 895 
0 1068 6 1 2 654 896 
0 1119 6 1 2 723 988 
0 1120 6 1 2 720 989 
0 1121 6 1 2 729 991 
0 1122 6 1 2 726 992 
0 1128 6 1 2 741 1002 
0 1129 6 1 2 738 1003 
0 1130 6 1 2 747 1005 
0 1131 6 1 2 744 1006 
0 1132 6 1 2 753 1008 
0 1133 6 1 2 750 1009 
0 1148 5 1 1 940 
0 1149 5 1 1 936 
0 1150 6 1 2 1054 1055 
0 1151 5 1 1 944 
0 1152 5 1 1 948 
0 1153 5 1 1 956 
0 1154 5 1 1 952 
0 1155 5 1 1 963 
0 1156 5 1 1 970 
0 1157 5 1 1 978 
0 1158 6 1 2 1063 1064 
0 1159 5 1 1 986 
0 1160 6 1 2 987 892 
0 1161 5 1 1 999 
0 1162 6 1 2 1067 1068 
0 1163 5 1 1 900 
0 1164 0 2 1 901 
2 1165 1 1164  
2 1166 1 1164  
0 1167 5 1 1 904 
0 1168 0 2 1 905 
2 1169 1 1168  
2 1170 1 1168  
0 1171 6 16 2 921 924 
2 1172 1 1171  
2 1173 1 1171  
2 1174 1 1171  
2 1175 1 1171  
2 1176 1 1171  
2 1177 1 1171  
2 1178 1 1171  
2 1179 1 1171  
2 1180 1 1171  
2 1181 1 1171  
2 1182 1 1171  
2 1183 1 1171  
2 1184 1 1171  
2 1185 1 1171  
2 1186 1 1171  
2 1187 1 1171  
0 1188 6 16 2 922 925 
2 1189 1 1188  
2 1190 1 1188  
2 1191 1 1188  
2 1192 1 1188  
2 1193 1 1188  
2 1194 1 1188  
2 1195 1 1188  
2 1196 1 1188  
2 1197 1 1188  
2 1198 1 1188  
2 1199 1 1188  
2 1200 1 1188  
2 1201 1 1188  
2 1202 1 1188  
2 1203 1 1188  
2 1204 1 1188  
0 1205 5 1 1 1011 
0 1206 6 1 2 1012 938 
0 1207 5 1 1 1014 
0 1208 6 1 2 1015 942 
0 1209 5 1 1 1017 
0 1210 6 1 2 1018 946 
0 1211 5 1 1 1020 
0 1212 6 1 2 1021 950 
0 1213 5 1 1 1023 
0 1214 6 1 2 1024 954 
0 1215 5 1 1 1026 
0 1216 6 1 2 1027 958 
0 1217 5 1 1 1029 
0 1218 5 1 1 960 
0 1219 5 1 1 1032 
0 1220 5 1 1 1035 
0 1221 6 1 2 1036 968 
0 1222 5 1 1 966 
0 1223 5 1 1 1038 
0 1224 6 1 2 1039 972 
0 1225 5 1 1 1041 
0 1226 6 1 2 1042 976 
0 1227 5 1 1 974 
0 1228 5 1 1 1044 
0 1229 6 1 2 1045 980 
0 1230 5 1 1 982 
0 1231 6 1 2 983 984 
0 1232 6 2 2 1119 1120 
2 1233 1 1232  
2 1234 1 1232  
0 1235 6 2 2 1121 1122 
2 1236 1 1235  
2 1237 1 1235  
0 1238 5 1 1 1047 
0 1239 6 1 2 1048 997 
0 1240 5 1 1 995 
0 1241 5 1 1 1050 
0 1242 6 1 2 1051 1001 
0 1243 6 2 2 1128 1129 
2 1244 1 1243  
2 1245 1 1243  
0 1246 6 2 2 1130 1131 
2 1247 1 1246  
2 1248 1 1246  
0 1249 6 2 2 1132 1133 
2 1250 1 1249  
2 1251 1 1249  
0 1252 0 2 1 908 
2 1253 1 1252  
2 1254 1 1252  
0 1255 0 2 1 909 
2 1256 1 1255  
2 1257 1 1255  
0 1258 0 2 1 911 
2 1259 1 1258  
2 1260 1 1258  
0 1261 0 2 1 912 
2 1262 1 1261  
2 1263 1 1261  
0 1264 5 2 1 1150 
2 1265 1 1264  
2 1266 1 1264  
0 1267 6 1 2 633 1159 
0 1309 6 1 2 690 1205 
0 1310 6 1 2 693 1207 
0 1311 6 1 2 696 1209 
0 1312 6 1 2 699 1211 
0 1313 6 1 2 702 1213 
0 1314 6 1 2 705 1215 
0 1315 6 1 2 708 1220 
0 1316 6 1 2 711 1223 
0 1317 6 1 2 714 1225 
0 1318 6 1 2 717 1228 
0 1319 5 2 1 1158 
2 1320 1 1319  
2 1321 1 1319  
0 1322 6 1 2 630 1230 
0 1327 6 1 2 732 1238 
0 1328 6 1 2 735 1241 
0 1334 5 2 1 1162 
2 1335 1 1334  
2 1336 1 1334  
0 1344 6 1 2 1267 1160 
0 1345 6 1 2 1250 894 
0 1346 5 1 1 1251 
0 1348 5 1 1 1256 
0 1349 5 1 1 1253 
0 1350 5 1 1 1262 
0 1351 5 1 1 1259 
0 1352 6 2 2 1309 1206 
2 1353 1 1352  
2 1354 1 1352  
0 1355 6 2 2 1310 1208 
2 1356 1 1355  
2 1357 1 1355  
0 1358 6 2 2 1311 1210 
2 1359 1 1358  
2 1360 1 1358  
0 1361 6 2 2 1312 1212 
2 1362 1 1361  
2 1363 1 1361  
0 1364 6 2 2 1313 1214 
2 1365 1 1364  
2 1366 1 1364  
0 1367 6 2 2 1314 1216 
2 1368 1 1367  
2 1369 1 1367  
0 1370 6 2 2 1315 1221 
2 1371 1 1370  
2 1372 1 1370  
0 1373 6 2 2 1316 1224 
2 1374 1 1373  
2 1375 1 1373  
0 1376 6 2 2 1317 1226 
2 1377 1 1376  
2 1378 1 1376  
0 1379 6 2 2 1318 1229 
2 1380 1 1379  
2 1381 1 1379  
0 1383 6 2 2 1322 1231 
2 1384 1 1383  
2 1385 1 1383  
0 1386 5 1 1 1233 
0 1387 6 1 2 1234 990 
0 1388 5 1 1 1236 
0 1389 6 1 2 1237 993 
0 1390 6 2 2 1327 1239 
2 1391 1 1390  
2 1392 1 1390  
0 1393 6 2 2 1328 1242 
2 1394 1 1393  
2 1395 1 1393  
0 1396 5 1 1 1244 
0 1397 6 1 2 1245 1004 
0 1398 5 1 1 1247 
0 1399 6 1 2 1248 1007 
0 1409 5 1 1 1320 
0 1412 6 1 2 651 1346 
0 1413 5 1 1 1335 
0 1416 0 2 1 1265 
2 1417 1 1416  
2 1418 1 1416  
0 1419 0 2 1 1266 
2 1420 1 1419  
2 1421 1 1419  
0 1433 6 1 2 636 1386 
0 1434 6 1 2 639 1388 
0 1438 6 1 2 642 1396 
0 1439 6 1 2 648 1398 
0 1440 5 2 1 1344 
2 1441 1 1440  
2 1442 1 1440  
0 1443 6 1 2 1356 1148 
0 1444 5 1 1 1357 
0 1445 6 1 2 1353 1149 
0 1446 5 1 1 1354 
0 1447 6 1 2 1359 1151 
0 1448 5 1 1 1360 
0 1451 6 1 2 1362 1152 
0 1452 5 1 1 1363 
0 1453 6 1 2 1368 1153 
0 1454 5 1 1 1369 
0 1455 6 1 2 1365 1154 
0 1456 5 1 1 1366 
0 1457 6 1 2 1374 1156 
0 1458 5 1 1 1375 
0 1459 6 1 2 1380 1157 
0 1460 5 1 1 1381 
0 1461 5 1 1 1384 
0 1462 6 1 2 1394 1161 
0 1463 5 1 1 1395 
0 1464 6 1 2 1345 1412 
0 1468 5 1 1 1371 
0 1469 6 1 2 1372 1222 
0 1470 5 1 1 1377 
0 1471 6 1 2 1378 1227 
0 1472 6 2 2 1387 1433 
2 1473 1 1472  
2 1474 1 1472  
0 1475 5 1 1 1391 
0 1476 6 1 2 1392 1240 
0 1478 6 2 2 1389 1434 
2 1479 1 1478  
2 1480 1 1478  
0 1481 6 2 2 1399 1439 
2 1482 1 1481  
2 1483 1 1481  
0 1484 6 2 2 1397 1438 
2 1485 1 1484  
2 1486 1 1484  
0 1487 6 1 2 941 1444 
0 1488 6 1 2 937 1446 
0 1489 6 1 2 945 1448 
0 1490 5 1 1 1420 
0 1491 5 1 1 1417 
0 1492 6 1 2 949 1452 
0 1493 6 1 2 957 1454 
0 1494 6 1 2 953 1456 
0 1495 6 1 2 971 1458 
0 1496 6 1 2 979 1460 
0 2739 6 1 2 2662 546 
0 1498 6 1 2 1000 1463 
0 1499 5 1 1 1441 
0 1500 6 1 2 967 1468 
0 1501 6 1 2 975 1470 
0 1504 6 1 2 996 1475 
0 2742 5 1 1 2666 
0 1510 5 2 1 1464 
2 1511 1 1510  
2 1512 1 1510  
0 1513 6 1 2 1443 1487 
0 1514 6 2 2 1445 1488 
2 1515 1 1514  
2 1516 1 1514  
0 1517 6 2 2 1447 1489 
2 1518 1 1517  
2 1519 1 1517  
0 1520 6 1 2 1451 1492 
0 1521 6 1 2 1453 1493 
0 1522 6 3 2 1455 1494 
2 1523 1 1522  
2 1524 1 1522  
2 1525 1 1522  
0 2745 6 1 8 2538 2541 2544 2547 2595 2598 2601 2604 
0 1526 6 1 2 1457 1495 
0 1527 6 1 2 1459 1496 
0 1528 5 1 1 1473 
0 1529 6 1 2 1462 1498 
0 1530 5 1 1 1479 
0 1531 5 1 1 1482 
0 1532 5 1 1 1485 
0 1534 6 2 2 1471 1501 
2 1535 1 1534  
2 1536 1 1534  
0 1537 6 2 2 1469 1500 
2 1538 1 1537  
2 1539 1 1537  
0 1540 6 2 2 1476 1504 
2 1541 1 1540  
2 1542 1 1540  
0 1546 5 2 1 1513 
2 1547 1 1546  
2 1548 1 1546  
0 1554 5 2 1 1521 
2 1555 1 1554  
2 1556 1 1554  
0 1557 5 3 1 1526 
2 1558 1 1557  
2 1559 1 1557  
2 1560 1 1557  
0 1561 5 2 1 1520 
2 1562 1 1561  
2 1563 1 1561  
0 1567 6 1 2 1486 1531 
0 1568 6 1 2 1483 1532 
0 1569 5 1 1 1511 
0 1571 5 2 1 1527 
2 1572 1 1571  
2 1573 1 1571  
0 1576 5 2 1 1529 
2 1577 1 1576  
2 1578 1 1576  
0 1588 0 2 1 1523 
2 1589 1 1588  
2 1590 1 1588  
0 1591 5 1 1 1535 
0 1593 5 1 1 1538 
0 1594 6 1 2 1541 1530 
0 1595 5 1 1 1542 
0 1596 6 2 2 1567 1568 
2 1597 1 1596  
2 1598 1 1596  
0 2760 6 1 2 366 2731 
0 1600 0 2 1 1518 
2 1601 1 1600  
2 1602 1 1600  
0 1603 0 2 1 1519 
2 1604 1 1603  
2 1605 1 1603  
0 1606 0 2 1 1524 
2 1607 1 1606  
2 1608 1 1606  
0 1609 0 2 1 1525 
2 1610 1 1609  
2 1611 1 1609  
0 1612 0 2 1 1515 
2 1613 1 1612  
2 1614 1 1612  
0 2763 6 1 2 375 2736 
0 1615 0 2 1 1516 
2 1616 1 1615  
2 1617 1 1615  
0 1620 0 2 1 1558 
2 1621 1 1620  
2 1622 1 1620  
0 1623 0 2 1 1555 
2 1624 1 1623  
2 1625 1 1623  
0 2766 6 1 2 384 2742 
0 1635 5 1 1 1572 
0 1636 6 1 2 1480 1595 
0 1638 6 1 2 1577 1569 
0 1639 5 1 1 1578 
0 1640 0 2 1 1562 
2 1641 1 1640  
2 1642 1 1640  
0 1643 0 2 1 1563 
2 1644 1 1643  
2 1645 1 1643  
0 1647 0 2 1 1547 
2 1648 1 1647  
2 1649 1 1647  
0 1651 0 2 1 1548 
2 1652 1 1651  
2 1653 1 1651  
0 1658 0 2 1 1556 
2 1659 1 1658  
2 1660 1 1658  
0 1661 0 2 1 1559 
2 1662 1 1661  
2 1663 1 1661  
0 1664 0 2 1 1560 
2 1665 1 1664  
2 1666 1 1664  
0 1671 6 1 2 1597 893 
0 1672 5 1 1 1598 
0 1675 5 1 1 1601 
0 1677 5 1 1 1604 
0 1678 6 1 2 1607 1217 
0 1679 5 1 1 1608 
0 1680 6 1 2 1610 1219 
0 1681 5 1 1 1611 
0 1682 5 1 1 1613 
0 1683 5 1 1 1616 
0 1685 6 2 2 1594 1636 
2 1686 1 1685  
2 1687 1 1685  
0 1688 6 1 2 1512 1639 
0 1697 0 2 1 1589 
2 1698 1 1697  
2 1699 1 1697  
0 1701 0 2 1 1590 
2 1702 1 1701  
2 1703 1 1701  
0 1706 6 1 2 645 1672 
0 1707 5 1 1 1644 
0 1708 6 1 2 1648 1675 
0 1709 5 1 1 1649 
0 1710 6 1 2 1652 1677 
0 1711 5 1 1 1653 
0 1712 6 1 2 1030 1679 
0 1713 6 1 2 1033 1681 
0 1714 0 2 1 1621 
2 1715 1 1714  
2 1716 1 1714  
0 1717 0 2 1 1622 
2 1718 1 1717  
2 1719 1 1717  
0 1720 6 1 2 1659 1593 
0 1721 5 1 1 1660 
0 1723 6 2 2 1638 1688 
2 1724 1 1723  
2 1725 1 1723  
0 1727 5 1 1 1662 
0 1728 5 1 1 1641 
0 1730 5 1 1 1665 
0 1731 0 2 1 1624 
2 1732 1 1731  
2 1733 1 1731  
0 1734 0 2 1 1625 
2 1735 1 1734  
2 1736 1 1734  
0 1740 6 1 2 1686 1528 
0 1741 5 1 1 1687 
0 1742 6 2 2 1671 1706 
2 1743 1 1742  
2 1744 1 1742  
0 1746 6 1 2 1602 1709 
0 1747 6 1 2 1605 1711 
0 1748 6 2 2 1678 1712 
2 1749 1 1748  
2 1750 1 1748  
0 1751 6 2 2 1680 1713 
2 1752 1 1751  
2 1753 1 1751  
0 1759 6 1 2 1539 1721 
0 1761 5 1 1 1698 
0 1762 6 1 2 1699 1727 
0 1763 5 1 1 1702 
0 1764 6 1 2 1703 1730 
0 1768 5 1 1 1718 
0 1769 6 1 2 1474 1741 
0 1772 6 1 2 1724 1413 
0 1773 5 1 1 1725 
0 1774 6 2 2 1708 1746 
2 1775 1 1774  
2 1776 1 1774  
0 1777 6 2 2 1710 1747 
2 1778 1 1777  
2 1779 1 1777  
0 1783 5 1 1 1732 
0 1784 6 1 2 1733 1682 
0 1785 5 1 1 1715 
0 1786 5 1 1 1735 
0 1787 6 1 2 1736 1683 
0 1788 6 2 2 1720 1759 
2 1789 1 1788  
2 1790 1 1788  
0 1791 6 1 2 1663 1761 
0 1792 6 1 2 1666 1763 
0 1795 6 1 2 1752 1155 
0 1796 5 1 1 1753 
0 1798 6 2 2 1740 1769 
2 1799 1 1798  
2 1800 1 1798  
0 1801 6 1 2 1336 1773 
0 1802 6 2 2 1743 291 
2 1803 1 1802  
2 1804 1 1802  
0 1807 5 1 1 1749 
0 1808 6 1 2 1750 1218 
0 1809 6 1 2 1614 1783 
0 1810 6 1 2 1617 1786 
0 1812 6 2 2 1791 1762 
2 1813 1 1812  
2 1814 1 1812  
0 1815 6 2 2 1792 1764 
2 1816 1 1815  
2 1817 1 1815  
0 1818 0 2 1 1744 
2 1819 1 1818  
2 1820 1 1818  
0 1821 6 1 2 1778 1490 
0 1822 5 1 1 1779 
0 1823 6 1 2 1775 1491 
0 1824 5 1 1 1776 
0 1825 6 1 2 964 1796 
0 1826 6 1 2 1789 1409 
0 1827 5 1 1 1790 
0 1830 6 2 2 1772 1801 
2 1831 1 1830  
2 1832 1 1830  
0 1837 6 1 2 961 1807 
0 1838 6 2 2 1809 1784 
2 1839 1 1838  
2 1840 1 1838  
0 1841 6 2 2 1810 1787 
2 1842 1 1841  
2 1843 1 1841  
0 1848 6 1 2 1421 1822 
0 1849 6 1 2 1418 1824 
0 1850 6 1 2 1795 1825 
0 1852 6 1 2 1321 1827 
0 1855 6 1 2 1816 1707 
0 1856 5 1 1 1817 
0 1857 5 1 1 1819 
0 1858 6 2 2 1799 292 
2 1859 1 1858  
2 1860 1 1858  
0 1864 5 1 1 1813 
0 1865 6 1 2 1814 1728 
0 1866 0 2 1 1800 
2 1867 1 1866  
2 1868 1 1866  
0 1869 0 2 1 1803 
2 1870 1 1869  
2 1871 1 1869  
0 1872 0 2 1 1804 
2 1873 1 1872  
2 1874 1 1872  
0 1875 6 2 2 1808 1837 
2 1876 1 1875  
2 1877 1 1875  
0 1878 6 1 2 1821 1848 
0 1879 6 2 2 1823 1849 
2 1880 1 1879  
2 1881 1 1879  
0 1882 6 1 2 1842 1768 
0 1883 5 1 1 1843 
0 1884 6 1 2 1826 1852 
0 1885 6 1 2 1645 1856 
0 1889 6 2 2 1831 293 
2 1890 1 1889  
2 1891 1 1889  
0 1895 5 1 1 1839 
0 1896 6 1 2 1840 1785 
0 1897 6 1 2 1642 1864 
0 1898 5 2 1 1850 
2 1899 1 1898  
2 1900 1 1898  
0 1902 0 2 1 1832 
2 1903 1 1902  
2 1904 1 1902  
0 1910 5 1 1 1878 
0 1911 6 1 2 1719 1883 
0 1912 5 1 1 1884 
0 1913 6 1 2 1855 1885 
0 1915 5 1 1 1867 
0 1919 6 1 2 1873 919 
0 1920 5 1 1 1874 
0 1921 6 1 2 1870 920 
0 1922 5 1 1 1871 
0 1923 5 1 1 1876 
0 1924 6 1 2 1716 1895 
0 1927 0 2 1 1859 
2 1928 1 1927  
2 1929 1 1927  
0 1930 0 2 1 1860 
2 1931 1 1930  
2 1932 1 1930  
0 1933 6 2 2 1865 1897 
2 1934 1 1933  
2 1935 1 1933  
0 1936 6 1 2 1882 1911 
0 1937 5 1 1 1899 
0 1938 5 1 1 1903 
0 1941 6 1 2 681 1920 
0 1942 6 1 2 678 1922 
0 1944 0 2 1 1880 
2 1945 1 1944  
2 1946 1 1944  
0 1947 5 2 1 1913 
2 1948 1 1947  
2 1949 1 1947  
0 1950 0 2 1 1890 
2 1951 1 1950  
2 1952 1 1950  
0 1953 0 2 1 1891 
2 1954 1 1953  
2 1955 1 1953  
0 1958 0 2 1 1881 
2 1959 1 1958  
2 1960 1 1958  
0 1961 6 2 2 1896 1924 
2 1962 1 1961  
2 1963 1 1961  
0 1965 7 2 2 1910 601 
2 1966 1 1965  
2 1967 1 1965  
0 1968 7 2 2 602 1912 
2 1969 1 1968  
2 1970 1 1968  
0 1975 6 1 2 1931 917 
0 1976 5 1 1 1932 
0 1977 6 1 2 1928 918 
0 1978 5 1 1 1929 
0 1979 6 1 2 1919 1941 
0 1980 6 2 2 1921 1942 
2 1981 1 1980  
2 1982 1 1980  
0 1985 5 1 1 1934 
0 1987 5 2 1 1936 
2 1988 1 1987  
2 1989 1 1987  
0 1999 5 1 1 1945 
0 2000 6 1 2 1946 1937 
0 2002 5 1 1 1948 
0 2003 6 1 2 1949 1499 
0 2004 6 1 2 1954 1350 
0 2005 5 1 1 1955 
0 2006 6 1 2 1951 1351 
0 2007 5 1 1 1952 
0 2008 6 1 2 675 1976 
0 2009 6 1 2 672 1978 
0 2012 5 1 1 1979 
0 2013 5 1 1 1959 
0 2014 6 1 2 1960 1923 
0 2015 5 1 1 1962 
0 2016 6 1 2 1963 1635 
0 2018 5 1 1 1966 
0 2019 5 1 1 1969 
0 2020 6 1 2 1900 1999 
0 2021 5 1 1 1988 
0 2022 6 1 2 1989 1591 
0 2023 6 1 2 1442 2002 
0 2024 6 1 2 1263 2005 
0 2025 6 1 2 1260 2007 
0 2026 6 1 2 1975 2008 
0 2027 6 2 2 1977 2009 
2 2028 1 2027  
2 2029 1 2027  
0 2030 5 2 1 1981 
2 2031 1 2030  
2 2032 1 2030  
0 2033 0 2 1 1982 
2 2034 1 2033  
2 2035 1 2033  
0 2036 6 1 2 1877 2013 
0 2037 6 1 2 1573 2015 
0 2038 6 1 2 2020 2000 
0 2039 6 1 2 1536 2021 
0 2040 6 1 2 2023 2003 
0 2041 6 1 2 2004 2024 
0 2042 6 2 2 2006 2025 
2 2043 1 2042  
2 2044 1 2042  
0 2047 5 1 1 2026 
