1	1	0	3	0	
1	5	0	3	0	
1	9	0	3	0	
1	13	0	3	0	
1	17	0	3	0	
1	21	0	3	0	
1	25	0	3	0	
1	29	0	3	0	
1	33	0	3	0	
1	37	0	3	0	
1	41	0	3	0	
1	45	0	3	0	
1	49	0	3	0	
1	53	0	3	0	
1	57	0	3	0	
1	61	0	3	0	
1	65	0	3	0	
1	69	0	3	0	
1	73	0	3	0	
1	77	0	3	0	
1	81	0	3	0	
1	85	0	3	0	
1	89	0	3	0	
1	93	0	3	0	
1	97	0	3	0	
1	101	0	3	0	
1	105	0	3	0	
1	109	0	3	0	
1	113	0	3	0	
1	117	0	3	0	
1	121	0	3	0	
1	125	0	3	0	
1	129	0	1	0	
1	130	0	1	0	
1	131	0	1	0	
1	132	0	1	0	
1	133	0	1	0	
1	134	0	1	0	
1	135	0	1	0	
1	136	0	1	0	
1	137	0	8	0	
0	250	2	1	2	756	759	
0	251	2	1	2	762	765	
0	252	2	1	2	768	771	
0	253	2	1	2	774	777	
0	254	2	1	2	780	783	
0	255	2	1	2	786	789	
0	256	2	1	2	792	795	
0	257	2	1	2	798	801	
0	258	2	1	2	804	807	
0	259	2	1	2	810	813	
0	260	2	1	2	816	819	
0	261	2	1	2	822	825	
0	262	2	1	2	828	839	
0	263	2	1	2	842	849	
0	264	2	1	2	852	859	
0	265	2	1	2	866	873	
0	266	7	1	2	129	880	
0	267	7	1	2	130	881	
0	268	7	1	2	131	882	
0	269	7	1	2	132	883	
0	270	7	1	2	133	884	
0	271	7	1	2	134	885	
0	272	7	1	2	135	886	
0	273	7	1	2	136	887	
0	274	2	1	2	757	769	
0	275	2	1	2	781	793	
0	276	2	1	2	760	772	
0	277	2	1	2	784	796	
0	278	2	1	2	763	775	
0	279	2	1	2	787	799	
0	280	2	1	2	766	778	
0	281	2	1	2	790	802	
0	282	2	1	2	805	817	
0	283	2	1	2	829	853	
0	284	2	1	2	808	820	
0	285	2	1	2	840	860	
0	286	2	1	2	811	823	
0	287	2	1	2	843	867	
0	288	2	1	2	814	826	
0	289	2	1	2	850	874	
0	290	2	2	2	250	251	
0	293	2	2	2	252	253	
0	296	2	2	2	254	255	
0	299	2	2	2	256	257	
0	302	2	2	2	258	259	
0	305	2	2	2	260	261	
0	308	2	2	2	262	263	
0	311	2	2	2	264	265	
0	314	2	1	2	274	275	
0	315	2	1	2	276	277	
0	316	2	1	2	278	279	
0	317	2	1	2	280	281	
0	318	2	1	2	282	283	
0	319	2	1	2	284	285	
0	320	2	1	2	286	287	
0	321	2	1	2	288	289	
0	338	2	1	2	900	902	
0	339	2	1	2	904	906	
0	340	2	1	2	901	905	
0	341	2	1	2	903	907	
0	342	2	1	2	908	910	
0	343	2	1	2	912	914	
0	344	2	1	2	909	913	
0	345	2	1	2	911	915	
0	346	2	1	2	266	342	
0	347	2	1	2	267	343	
0	348	2	1	2	268	344	
0	349	2	1	2	269	345	
0	350	2	1	2	270	338	
0	351	2	1	2	271	339	
0	352	2	1	2	272	340	
0	353	2	1	2	273	341	
0	354	2	12	2	314	346	
0	367	2	12	2	315	347	
0	380	2	12	2	316	348	
0	393	2	12	2	317	349	
0	406	2	12	2	318	350	
0	419	2	12	2	319	351	
0	432	2	12	2	320	352	
0	445	2	12	2	321	353	
0	554	5	1	1	916	
0	555	5	1	1	928	
0	556	5	1	1	940	
0	557	5	1	1	917	
0	558	5	1	1	929	
0	559	5	1	1	952	
0	560	5	1	1	918	
0	561	5	1	1	941	
0	562	5	1	1	953	
0	563	5	1	1	930	
0	564	5	1	1	942	
0	565	5	1	1	954	
0	566	5	1	1	976	
0	567	5	1	1	1000	
0	568	5	1	1	977	
0	569	5	1	1	988	
0	570	5	1	1	964	
0	571	5	1	1	1001	
0	572	5	1	1	965	
0	573	5	1	1	989	
0	574	5	1	1	966	
0	575	5	1	1	978	
0	576	5	1	1	990	
0	577	5	1	1	967	
0	578	5	1	1	979	
0	579	5	1	1	1002	
0	580	5	1	1	968	
0	581	5	1	1	991	
0	582	5	1	1	1003	
0	583	5	1	1	980	
0	584	5	1	1	992	
0	585	5	1	1	1004	
0	586	5	1	1	931	
0	587	5	1	1	955	
0	588	5	1	1	932	
0	589	5	1	1	943	
0	590	5	1	1	919	
0	591	5	1	1	956	
0	592	5	1	1	920	
0	593	5	1	1	944	
0	594	7	1	4	554	555	556	957	
0	595	7	1	4	557	558	945	559	
0	596	7	1	4	560	933	561	562	
0	597	7	1	4	921	563	564	565	
0	598	7	1	4	574	575	576	1005	
0	599	7	1	4	577	578	993	579	
0	600	7	1	4	580	981	581	582	
0	601	7	1	4	969	583	584	585	
0	602	3	4	4	594	595	596	597	
0	607	3	4	4	598	599	600	601	
0	620	7	4	5	970	566	994	567	831	
0	625	7	4	5	971	568	569	1006	832	
0	630	7	4	5	570	982	995	571	833	
0	635	7	4	5	572	983	573	1007	834	
0	640	7	4	5	922	586	946	587	835	
0	645	7	4	5	923	588	589	958	836	
0	650	7	4	5	590	934	947	591	837	
0	655	7	4	5	592	935	593	959	838	
0	692	7	1	2	924	845	
0	693	7	1	2	936	846	
0	694	7	1	2	948	847	
0	695	7	1	2	960	848	
0	696	7	1	2	925	855	
0	697	7	1	2	937	856	
0	698	7	1	2	949	857	
0	699	7	1	2	961	858	
0	700	7	1	2	926	862	
0	701	7	1	2	938	863	
0	702	7	1	2	950	864	
0	703	7	1	2	962	865	
0	704	7	1	2	927	869	
0	705	7	1	2	939	870	
0	706	7	1	2	951	871	
0	707	7	1	2	963	872	
0	708	7	1	2	972	876	
0	709	7	1	2	984	877	
0	710	7	1	2	996	878	
0	711	7	1	2	1008	879	
0	712	7	1	2	973	888	
0	713	7	1	2	985	889	
0	714	7	1	2	997	890	
0	715	7	1	2	1009	891	
0	716	7	1	2	974	892	
0	717	7	1	2	986	893	
0	718	7	1	2	998	894	
0	719	7	1	2	1010	895	
0	720	7	1	2	975	896	
0	721	7	1	2	987	897	
0	722	7	1	2	999	898	
0	723	7	1	2	1011	899	
3	724	2	0	2	758	692	
3	725	2	0	2	761	693	
3	726	2	0	2	764	694	
3	727	2	0	2	767	695	
3	728	2	0	2	770	696	
3	729	2	0	2	773	697	
3	730	2	0	2	776	698	
3	731	2	0	2	779	699	
3	732	2	0	2	782	700	
3	733	2	0	2	785	701	
3	734	2	0	2	788	702	
3	735	2	0	2	791	703	
3	736	2	0	2	794	704	
3	737	2	0	2	797	705	
3	738	2	0	2	800	706	
3	739	2	0	2	803	707	
3	740	2	0	2	806	708	
3	741	2	0	2	809	709	
3	742	2	0	2	812	710	
3	743	2	0	2	815	711	
3	744	2	0	2	818	712	
3	745	2	0	2	821	713	
3	746	2	0	2	824	714	
3	747	2	0	2	827	715	
3	748	2	0	2	830	716	
3	749	2	0	2	841	717	
3	750	2	0	2	844	718	
3	751	2	0	2	851	719	
3	752	2	0	2	854	720	
3	753	2	0	2	861	721	
3	754	2	0	2	868	722	
3	755	2	0	2	875	723	
2	756	1	1			
2	757	1	1			
2	758	1	1			
2	759	1	5			
2	760	1	5			
2	761	1	5			
2	762	1	9			
2	763	1	9			
2	764	1	9			
2	765	1	13			
2	766	1	13			
2	767	1	13			
2	768	1	17			
2	769	1	17			
2	770	1	17			
2	771	1	21			
2	772	1	21			
2	773	1	21			
2	774	1	25			
2	775	1	25			
2	776	1	25			
2	777	1	29			
2	778	1	29			
2	779	1	29			
2	780	1	33			
2	781	1	33			
2	782	1	33			
2	783	1	37			
2	784	1	37			
2	785	1	37			
2	786	1	41			
2	787	1	41			
2	788	1	41			
2	789	1	45			
2	790	1	45			
2	791	1	45			
2	792	1	49			
2	793	1	49			
2	794	1	49			
2	795	1	53			
2	796	1	53			
2	797	1	53			
2	798	1	57			
2	799	1	57			
2	800	1	57			
2	801	1	61			
2	802	1	61			
2	803	1	61			
2	804	1	65			
2	805	1	65			
2	806	1	65			
2	807	1	69			
2	808	1	69			
2	809	1	69			
2	810	1	73			
2	811	1	73			
2	812	1	73			
2	813	1	77			
2	814	1	77			
2	815	1	77			
2	816	1	81			
2	817	1	81			
2	818	1	81			
2	819	1	85			
2	820	1	85			
2	821	1	85			
2	822	1	89			
2	823	1	89			
2	824	1	89			
2	825	1	93			
2	826	1	93			
2	827	1	93			
2	828	1	97			
2	829	1	97			
2	830	1	97			
2	831	1	602			
2	832	1	602			
2	833	1	602			
2	834	1	602			
2	835	1	607			
2	836	1	607			
2	837	1	607			
2	838	1	607			
2	839	1	101			
2	840	1	101			
2	841	1	101			
2	842	1	105			
2	843	1	105			
2	844	1	105			
2	845	1	620			
2	846	1	620			
2	847	1	620			
2	848	1	620			
2	849	1	109			
2	850	1	109			
2	851	1	109			
2	852	1	113			
2	853	1	113			
2	854	1	113			
2	855	1	625			
2	856	1	625			
2	857	1	625			
2	858	1	625			
2	859	1	117			
2	860	1	117			
2	861	1	117			
2	862	1	630			
2	863	1	630			
2	864	1	630			
2	865	1	630			
2	866	1	121			
2	867	1	121			
2	868	1	121			
2	869	1	635			
2	870	1	635			
2	871	1	635			
2	872	1	635			
2	873	1	125			
2	874	1	125			
2	875	1	125			
2	876	1	640			
2	877	1	640			
2	878	1	640			
2	879	1	640			
2	880	1	137			
2	881	1	137			
2	882	1	137			
2	883	1	137			
2	884	1	137			
2	885	1	137			
2	886	1	137			
2	887	1	137			
2	888	1	645			
2	889	1	645			
2	890	1	645			
2	891	1	645			
2	892	1	650			
2	893	1	650			
2	894	1	650			
2	895	1	650			
2	896	1	655			
2	897	1	655			
2	898	1	655			
2	899	1	655			
2	900	1	290			
2	901	1	290			
2	902	1	293			
2	903	1	293			
2	904	1	296			
2	905	1	296			
2	906	1	299			
2	907	1	299			
2	908	1	302			
2	909	1	302			
2	910	1	305			
2	911	1	305			
2	912	1	308			
2	913	1	308			
2	914	1	311			
2	915	1	311			
2	916	1	354			
2	917	1	354			
2	918	1	354			
2	919	1	354			
2	920	1	354			
2	921	1	354			
2	922	1	354			
2	923	1	354			
2	924	1	354			
2	925	1	354			
2	926	1	354			
2	927	1	354			
2	928	1	367			
2	929	1	367			
2	930	1	367			
2	931	1	367			
2	932	1	367			
2	933	1	367			
2	934	1	367			
2	935	1	367			
2	936	1	367			
2	937	1	367			
2	938	1	367			
2	939	1	367			
2	940	1	380			
2	941	1	380			
2	942	1	380			
2	943	1	380			
2	944	1	380			
2	945	1	380			
2	946	1	380			
2	947	1	380			
2	948	1	380			
2	949	1	380			
2	950	1	380			
2	951	1	380			
2	952	1	393			
2	953	1	393			
2	954	1	393			
2	955	1	393			
2	956	1	393			
2	957	1	393			
2	958	1	393			
2	959	1	393			
2	960	1	393			
2	961	1	393			
2	962	1	393			
2	963	1	393			
2	964	1	406			
2	965	1	406			
2	966	1	406			
2	967	1	406			
2	968	1	406			
2	969	1	406			
2	970	1	406			
2	971	1	406			
2	972	1	406			
2	973	1	406			
2	974	1	406			
2	975	1	406			
2	976	1	419			
2	977	1	419			
2	978	1	419			
2	979	1	419			
2	980	1	419			
2	981	1	419			
2	982	1	419			
2	983	1	419			
2	984	1	419			
2	985	1	419			
2	986	1	419			
2	987	1	419			
2	988	1	432			
2	989	1	432			
2	990	1	432			
2	991	1	432			
2	992	1	432			
2	993	1	432			
2	994	1	432			
2	995	1	432			
2	996	1	432			
2	997	1	432			
2	998	1	432			
2	999	1	432			
2	1000	1	445			
2	1001	1	445			
2	1002	1	445			
2	1003	1	445			
2	1004	1	445			
2	1005	1	445			
2	1006	1	445			
2	1007	1	445			
2	1008	1	445			
2	1009	1	445			
2	1010	1	445			
2	1011	1	445			
