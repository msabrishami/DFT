1	1	0	1	0	
1	2	0	1	0	
1	3	0	1	0	
1	4	0	1	0	
1	5	0	1	0	
1	6	0	1	0	
1	7	0	1	0	
1	8	0	16	0	
1	11	0	2	0	
1	14	0	1	0	
1	15	0	1	0	
1	16	0	11	0	
1	19	0	1	0	
1	20	0	1	0	
1	21	0	1	0	
1	22	0	1	0	
1	23	0	1	0	
1	24	0	1	0	
1	25	0	1	0	
1	26	0	1	0	
1	27	0	1	0	
1	28	0	1	0	
1	29	0	10	0	
1	32	0	1	0	
1	33	0	1	0	
1	34	0	1	0	
1	35	0	1	0	
1	36	0	1	0	
1	37	0	2	0	
1	40	0	2	0	
1	43	0	1	0	
1	44	0	2	0	
1	47	0	1	0	
1	48	0	1	0	
1	49	0	1	0	
1	50	0	1	0	
1	51	0	1	0	
1	52	0	1	0	
1	53	0	1	0	
1	54	0	1	0	
1	55	0	1	0	
1	56	0	1	0	
1	57	0	2	0	
1	60	0	1	0	
1	61	0	1	0	
1	62	0	1	0	
1	63	0	1	0	
1	64	0	1	0	
1	65	0	1	0	
1	66	0	1	0	
1	67	0	1	0	
1	68	0	1	0	
1	69	0	2	0	
1	72	0	1	0	
1	73	0	1	0	
1	74	0	1	0	
1	75	0	1	0	
1	76	0	1	0	
1	77	0	1	0	
1	78	0	1	0	
1	79	0	1	0	
1	80	0	1	0	
1	81	0	1	0	
1	82	0	2	0	
1	85	0	1	0	
1	86	0	1	0	
1	87	0	1	0	
1	88	0	1	0	
1	89	0	1	0	
1	90	0	1	0	
1	91	0	1	0	
1	92	0	1	0	
1	93	0	1	0	
1	94	0	1	0	
1	95	0	1	0	
1	96	0	2	0	
1	99	0	1	0	
1	100	0	1	0	
1	101	0	1	0	
1	102	0	1	0	
1	103	0	1	0	
1	104	0	1	0	
1	105	0	1	0	
1	106	0	1	0	
1	107	0	1	0	
1	108	0	2	0	
1	111	0	1	0	
1	112	0	1	0	
1	113	0	1	0	
1	114	0	1	0	
1	115	0	1	0	
1	116	0	1	0	
1	117	0	1	0	
1	118	0	1	0	
1	119	0	1	0	
1	120	0	2	0	
1	123	0	1	0	
1	124	0	1	0	
1	125	0	1	0	
1	126	0	1	0	
1	127	0	1	0	
1	128	0	1	0	
1	129	0	1	0	
1	130	0	1	0	
1	131	0	1	0	
1	132	0	2	0	
1	135	0	1	0	
1	136	0	1	0	
1	137	0	1	0	
1	138	0	1	0	
1	139	0	1	0	
1	140	0	1	0	
1	141	0	1	0	
1	142	0	1	0	
3	143	0	0	0	
3	144	0	0	0	
3	145	0	0	0	
3	146	0	0	0	
3	147	0	0	0	
3	148	0	0	0	
3	149	0	0	0	
3	150	0	0	0	
3	151	0	0	0	
3	152	0	0	0	
3	153	0	0	0	
3	154	0	0	0	
3	155	0	0	0	
3	156	0	0	0	
3	157	0	0	0	
3	158	0	0	0	
3	159	0	0	0	
3	160	0	0	0	
3	161	0	0	0	
3	162	0	0	0	
3	163	0	0	0	
3	164	0	0	0	
3	165	0	0	0	
3	166	0	0	0	
3	167	0	0	0	
3	168	0	0	0	
3	169	0	0	0	
3	170	0	0	0	
3	171	0	0	0	
3	172	0	0	0	
3	173	0	0	0	
3	174	0	0	0	
3	175	0	0	0	
3	176	0	0	0	
3	177	0	0	0	
3	178	0	0	0	
3	179	0	0	0	
3	180	0	0	0	
3	181	0	0	0	
3	182	0	0	0	
3	183	0	0	0	
3	184	0	0	0	
3	185	0	0	0	
3	186	0	0	0	
3	187	0	0	0	
3	188	0	0	0	
3	189	0	0	0	
3	190	0	0	0	
3	191	0	0	0	
3	192	0	0	0	
3	193	0	0	0	
3	194	0	0	0	
3	195	0	0	0	
3	196	0	0	0	
3	197	0	0	0	
3	198	0	0	0	
3	199	0	0	0	
3	200	0	0	0	
3	201	0	0	0	
3	202	0	0	0	
3	203	0	0	0	
3	204	0	0	0	
3	205	0	0	0	
3	206	0	0	0	
3	207	0	0	0	
3	208	0	0	0	
3	209	0	0	0	
3	210	0	0	0	
3	211	0	0	0	
3	212	0	0	0	
3	213	0	0	0	
3	214	0	0	0	
3	215	0	0	0	
3	216	0	0	0	
3	217	0	0	0	
3	218	0	0	0	
3	219	0	0	0	
1	224	0	2	0	
1	227	0	22	0	
1	230	0	1	0	
1	231	0	2	0	
1	234	0	22	0	
1	237	0	4	0	
1	241	0	4	0	
1	246	0	6	0	
3	253	0	0	0	
1	256	0	3	0	
1	259	0	3	0	
1	262	0	1	0	
1	263	0	3	0	
1	266	0	3	0	
1	269	0	3	0	
1	272	0	3	0	
1	275	0	3	0	
1	278	0	3	0	
1	281	0	3	0	
1	284	0	3	0	
1	287	0	3	0	
3	290	0	0	0	
1	294	0	3	0	
1	297	0	4	0	
1	301	0	4	0	
1	305	0	4	0	
1	309	0	4	0	
1	313	0	3	0	
1	316	0	3	0	
1	319	0	22	0	
1	322	0	22	0	
1	325	0	2	0	
1	328	0	2	0	
1	331	0	2	0	
1	334	0	2	0	
1	337	0	2	0	
1	340	0	2	0	
1	343	0	2	0	
1	346	0	2	0	
1	349	0	2	0	
1	352	0	2	0	
1	355	0	2	0	
0	405	7	1	2	1	3	
0	408	5	1	1	230	
0	425	5	1	1	262	
0	485	7	1	4	4129	4125	4119	4115	
0	486	5	1	1	405	
3	487	5	0	1	3944	
3	488	5	0	1	3985	
3	489	5	0	1	3965	
3	490	5	0	1	3967	
3	491	5	0	1	3952	
3	492	5	0	1	3983	
3	493	5	0	1	3946	
3	494	5	0	1	3977	
0	495	7	1	3	2	15	4061	
0	499	7	1	2	3938	3939	
0	533	5	3	1	4065	
0	537	5	5	1	4071	
0	543	7	1	2	3903	4072	
0	544	7	2	4	3986	3966	3968	3945	
0	547	7	2	4	3984	3947	3978	3953	
0	574	5	4	1	4079	
0	578	5	4	1	4082	
0	606	5	1	1	4213	
0	607	5	1	1	4215	
0	608	5	1	1	4221	
0	609	5	1	1	4223	
0	610	5	1	1	4225	
0	611	5	1	1	4227	
0	612	5	1	1	4239	
0	650	5	1	1	4241	
0	651	7	3	2	7	4062	
0	655	5	4	1	4085	
0	659	5	4	1	4088	
0	663	5	4	1	4091	
0	667	5	4	1	4094	
0	671	5	4	1	4097	
0	675	5	4	1	4100	
0	679	5	4	1	4103	
0	683	5	4	1	4106	
0	687	5	6	1	4109	
0	705	5	6	1	4112	
0	711	5	4	1	4116	
0	715	5	4	1	4120	
0	719	5	4	1	4126	
0	723	5	4	1	4130	
0	727	5	2	1	4161	
0	730	5	2	1	4164	
0	733	5	1	1	4229	
0	734	5	1	1	4237	
3	792	5	0	1	485	
3	799	5	0	1	495	
0	800	5	2	1	499	
0	900	6	1	2	4216	606	
0	901	6	1	2	4214	607	
0	902	6	1	2	4224	608	
0	903	6	1	2	4222	609	
0	904	6	1	2	4228	610	
0	905	6	1	2	4226	611	
0	998	6	1	2	4238	733	
0	999	6	1	2	4230	734	
3	1026	7	0	2	94	219	
0	1027	7	1	2	4211	4337	
3	1028	5	0	1	4338	
3	1029	6	0	2	4037	4339	
0	1032	5	1	1	4301	
0	1033	5	1	1	4303	
3	1034	7	0	2	4304	4302	
0	1042	5	10	1	4015	
0	1053	5	10	1	4039	
0	1064	7	1	3	80	4016	4040	
0	1065	7	1	3	68	4017	4041	
0	1066	7	1	3	79	4018	4042	
0	1067	7	1	3	78	4019	4043	
0	1068	7	1	3	77	4020	4044	
0	1069	7	1	2	3904	4296	
0	1075	5	10	1	4021	
0	1086	5	10	1	4045	
0	1097	7	1	3	76	4022	4046	
0	1098	7	1	3	75	4023	4047	
0	1099	7	1	3	74	4024	4048	
0	1100	7	1	3	73	4025	4049	
0	1101	7	1	3	72	4026	4050	
0	1102	5	10	1	4167	
0	1113	5	10	1	4189	
0	1124	7	1	3	114	4168	4190	
0	1125	7	1	3	113	4169	4191	
0	1126	7	1	3	112	4170	4192	
0	1127	7	1	3	111	4171	4193	
0	1128	7	1	2	4172	4194	
0	1129	6	3	2	900	901	
0	1133	6	3	2	902	903	
0	1137	6	4	2	904	905	
0	1140	5	1	1	4086	
0	1141	6	1	2	4087	612	
0	1142	5	1	1	4092	
0	1143	5	1	1	4089	
0	1144	5	1	1	4098	
0	1145	5	1	1	4095	
0	1146	5	10	1	4173	
0	1157	5	10	1	4195	
0	1168	7	1	3	118	4174	4196	
0	1169	7	1	3	107	4175	4197	
0	1170	7	1	3	117	4176	4198	
0	1171	7	1	3	116	4177	4199	
0	1172	7	1	3	115	4178	4200	
0	1173	5	4	1	3909	
0	1178	5	5	1	3910	
0	1184	5	1	1	4113	
0	1185	6	1	2	4114	650	
0	1186	5	1	1	4121	
0	1187	5	1	1	4117	
0	1188	5	1	1	4131	
0	1189	5	1	1	4127	
0	1200	5	4	1	3924	
0	1205	5	4	1	3925	
0	1210	5	1	1	4083	
0	1211	5	1	1	4080	
0	1212	5	1	1	4104	
0	1213	5	1	1	4101	
0	1214	5	1	1	4110	
0	1215	5	1	1	4107	
0	1216	6	2	2	998	999	
0	1249	5	1	1	4165	
0	1250	5	1	1	4162	
3	1269	5	0	1	1027	
0	1275	7	1	2	4212	1032	
0	1276	7	1	2	4038	1033	
0	1302	3	1	2	1069	543	
0	1351	6	1	2	4240	1140	
0	1352	6	1	2	4090	1142	
0	1353	6	1	2	4093	1143	
0	1354	6	1	2	4096	1144	
0	1355	6	1	2	4099	1145	
0	1395	6	1	2	4242	1184	
0	1396	6	1	2	4118	1186	
0	1397	6	1	2	4122	1187	
0	1398	6	1	2	4128	1188	
0	1399	6	1	2	4132	1189	
0	1422	6	1	2	4081	1210	
0	1423	6	1	2	4084	1211	
0	1424	6	1	2	4102	1212	
0	1425	6	1	2	4105	1213	
0	1426	6	1	2	4108	1214	
0	1427	6	1	2	4111	1215	
0	1440	6	1	2	4163	1249	
0	1441	6	1	2	4166	1250	
3	1448	5	0	1	1034	
0	1449	5	1	1	1275	
0	1450	5	1	1	1276	
0	1451	7	1	3	93	4494	4507	
0	1452	7	1	3	55	4027	4508	
0	1453	7	1	3	67	4495	4051	
0	1454	7	1	3	81	4496	4509	
0	1455	7	1	3	43	4028	4510	
0	1456	7	1	3	56	4497	4052	
0	1457	7	1	3	92	4498	4511	
0	1458	7	1	3	54	4029	4512	
0	1459	7	1	3	66	4499	4053	
0	1460	7	1	3	91	4500	4513	
0	1461	7	1	3	53	4030	4514	
0	1462	7	1	3	65	4501	4054	
0	1463	7	1	3	90	4502	4515	
0	1464	7	1	3	52	4031	4516	
0	1465	7	1	3	64	4503	4055	
0	1466	7	1	3	89	4525	4535	
0	1467	7	1	3	51	4032	4536	
0	1468	7	1	3	63	4526	4056	
0	1469	7	1	3	88	4527	4537	
0	1470	7	1	3	50	4033	4538	
0	1471	7	1	3	62	4528	4057	
0	1472	7	1	3	87	4529	4539	
0	1473	7	1	3	49	4034	4540	
0	1474	7	1	2	4530	4058	
0	1475	7	1	3	86	4531	4541	
0	1476	7	1	3	48	4035	4542	
0	1477	7	1	3	61	4532	4059	
0	1478	7	1	3	85	4533	4543	
0	1479	7	1	3	47	4036	4544	
0	1480	7	1	3	60	4534	4060	
0	1481	7	1	3	138	4554	4579	
0	1482	7	1	3	102	4179	4580	
0	1483	7	1	3	126	4555	4201	
0	1484	7	1	3	137	4556	4581	
0	1485	7	1	3	101	4180	4582	
0	1486	7	1	3	125	4557	4202	
0	1487	7	1	3	136	4558	4583	
0	1488	7	1	3	100	4181	4584	
0	1489	7	1	3	124	4559	4203	
0	1490	7	1	3	135	4560	4585	
0	1491	7	1	3	99	4182	4586	
0	1492	7	1	3	123	4561	4204	
0	1493	7	1	2	4562	4587	
0	1494	7	1	2	4183	4588	
0	1495	7	1	2	4563	4205	
0	1496	5	2	1	4598	
0	1499	5	2	1	4604	
0	1502	6	3	2	1351	1141	
0	1506	6	3	2	1352	1353	
0	1510	6	4	2	1354	1355	
0	1519	5	1	1	4314	
0	1520	5	1	1	4321	
0	1521	5	1	1	4340	
0	1522	5	1	1	4346	
0	1523	5	1	1	4350	
0	1524	5	1	1	4354	
0	1525	5	1	1	4358	
0	1526	5	1	1	4362	
0	1527	5	1	1	4366	
0	1528	5	1	1	4370	
0	1529	7	1	3	142	4613	4623	
0	1530	7	1	3	106	4184	4624	
0	1531	7	1	3	130	4614	4206	
0	1532	7	1	3	131	4615	4625	
0	1533	7	1	3	95	4185	4626	
0	1534	7	1	3	119	4616	4207	
0	1535	7	1	3	141	4617	4627	
0	1536	7	1	3	105	4186	4628	
0	1537	7	1	3	129	4618	4208	
0	1538	7	1	3	140	4619	4629	
0	1539	7	1	3	104	4187	4630	
0	1540	7	1	3	128	4620	4209	
0	1541	7	1	3	139	4621	4631	
0	1542	7	1	3	103	4188	4632	
0	1543	7	1	3	127	4622	4210	
0	1544	7	1	2	19	4633	
0	1545	7	1	2	4	4634	
0	1546	7	1	2	20	4635	
0	1547	7	1	2	5	4636	
0	1548	7	1	2	21	4637	
0	1549	7	1	2	22	4638	
0	1550	7	1	2	23	4639	
0	1551	7	1	2	6	4640	
0	1552	7	1	2	24	4641	
0	1553	6	3	2	1395	1185	
0	1557	6	3	2	1396	1397	
0	1561	6	4	2	1398	1399	
0	1564	7	1	2	25	4646	
0	1565	7	1	2	32	4647	
0	1566	7	1	2	26	4648	
0	1567	7	1	2	33	4649	
0	1568	7	1	2	27	4650	
0	1569	7	1	2	34	4651	
0	1570	7	1	2	35	4652	
0	1571	7	1	2	28	4653	
0	1572	5	1	1	4374	
0	1573	5	1	1	4380	
0	1574	5	1	1	4386	
0	1575	5	1	1	4390	
0	1576	5	1	1	4394	
0	1577	5	1	1	4398	
0	1578	6	2	2	1422	1423	
0	1581	5	1	1	4654	
0	1582	6	2	2	1426	1427	
0	1585	6	2	2	1424	1425	
0	1588	6	2	2	1440	1441	
3	1591	7	0	2	1449	1450	
0	1596	3	5	4	1451	1452	1453	1064	
0	1600	3	6	4	1454	1455	1456	1065	
0	1606	3	5	4	1457	1458	1459	1066	
3	1612	3	0	4	1460	1461	1462	1067	
3	1615	3	0	4	1463	1464	1465	1068	
3	1619	3	0	4	1466	1467	1468	1097	
3	1624	3	0	4	1469	1470	1471	1098	
3	1628	3	0	4	1472	1473	1474	1099	
3	1631	3	0	4	1475	1476	1477	1100	
3	1634	3	0	4	1478	1479	1480	1101	
0	1637	3	5	4	1481	1482	1483	1124	
0	1642	3	5	4	1484	1485	1486	1125	
0	1647	3	4	4	1487	1488	1489	1126	
0	1651	3	5	4	1490	1491	1492	1127	
0	1656	3	4	4	1493	1494	1495	1128	
0	1676	3	5	4	1532	1533	1534	1169	
0	1681	3	5	4	1535	1536	1537	1170	
0	1686	3	5	4	1538	1539	1540	1171	
0	1690	3	3	4	1541	1542	1543	1172	
0	1708	3	2	4	1529	1530	1531	1168	
0	1770	5	2	1	4692	
0	1773	5	2	1	4695	
0	1776	5	1	1	4609	
0	1777	5	1	1	4610	
0	1784	7	1	3	4605	4599	4611	
0	1785	7	1	3	4690	4688	4612	
0	1795	5	2	1	4702	
0	1798	5	2	1	4705	
0	1807	5	1	1	4726	
0	1808	5	1	1	4716	
0	1809	6	1	2	4717	1581	
0	1810	5	1	1	4718	
0	1811	5	1	1	4724	
0	1813	7	1	2	4738	4066	
0	1814	7	1	2	4756	4067	
0	1815	7	1	2	4745	4068	
3	1816	5	0	1	4804	
3	1817	5	0	1	4809	
3	1818	5	0	1	4799	
3	1819	5	0	1	4780	
3	1820	5	0	1	4772	
3	1821	5	0	1	4768	
0	1822	7	1	4	4063	4013	36	4728	
0	1823	7	1	4	4064	4014	4729	486	
0	1827	5	2	1	4757	
0	1830	7	1	2	4746	4297	
0	1831	7	1	2	4758	4298	
0	1832	7	1	2	4773	4073	
0	1833	5	4	1	4739	
0	1836	5	6	1	4747	
0	1841	5	10	1	4759	
0	1885	6	2	2	4402	4813	
0	1888	6	2	2	4404	4818	
0	1894	7	2	2	4800	425	
0	1897	5	2	1	4805	
0	1908	7	1	3	4689	4606	1776	
0	1909	7	1	3	4600	4691	1777	
0	1910	7	1	2	4748	3911	
0	1911	7	1	2	4760	3912	
0	1912	7	1	2	4765	3913	
0	1913	7	1	2	4769	3914	
0	1914	7	1	2	4774	3915	
0	1915	7	1	2	4781	3916	
0	1916	7	1	2	4787	3917	
0	1917	7	1	2	4791	3918	
0	1918	7	1	2	4795	3919	
0	1919	5	1	1	4847	
0	1928	7	1	2	4824	3926	
0	1929	7	1	2	4829	3927	
0	1930	7	1	2	4834	3928	
0	1931	7	1	2	4839	3929	
0	1932	7	1	2	4801	3930	
0	1933	7	1	2	4806	3931	
0	1934	7	1	2	4810	3932	
0	1935	7	1	2	4814	3933	
0	1939	6	1	2	4655	1808	
0	1940	6	1	2	4725	1810	
0	1941	6	1	2	4719	1811	
3	1969	3	0	2	4293	1815	
3	1970	5	0	1	1822	
3	1971	5	0	1	1823	
0	2028	5	1	1	4698	
0	2029	5	1	1	4699	
0	2030	4	1	2	1908	1784	
0	2031	4	1	2	1909	1785	
0	2032	7	1	3	4696	4693	4700	
0	2033	7	1	3	4865	4863	4701	
0	2034	3	1	2	1571	1935	
0	2040	5	1	1	4708	
0	2041	5	1	1	4709	
0	2042	7	1	3	4706	4703	4710	
0	2043	7	1	3	4879	4875	4711	
0	2046	6	2	2	1939	1809	
0	2049	6	2	2	1940	1941	
0	2052	3	2	2	1544	1910	
0	2055	3	2	2	1545	1911	
0	2058	3	2	2	1546	1912	
0	2061	3	2	2	1547	1913	
0	2064	3	2	2	1548	1914	
0	2067	3	2	2	1549	1915	
0	2070	3	2	2	1550	1916	
0	2073	3	2	2	1551	1917	
0	2076	3	2	2	1552	1918	
0	2079	3	2	2	1564	1928	
0	2095	3	2	2	1565	1929	
0	2098	3	2	2	1566	1930	
0	2101	3	2	2	1567	1931	
0	2104	3	2	2	1568	1932	
0	2107	3	2	2	1569	1933	
0	2110	3	2	2	1570	1934	
0	2113	7	9	3	4920	4918	3942	
0	2119	5	1	1	4919	
0	2120	6	6	2	408	4892	
0	2125	7	1	2	4740	4299	
0	2126	7	1	2	4770	4074	
0	2127	7	1	2	4766	4300	
0	2128	5	10	1	4767	
0	2135	5	8	1	4771	
0	2141	5	4	1	4782	
0	2144	5	4	1	4788	
0	2147	5	4	1	4792	
0	2150	5	4	1	4796	
0	2153	7	1	2	4403	4914	
0	2154	7	1	2	4915	4815	
0	2155	7	1	2	4405	4916	
0	2156	7	1	2	4917	4819	
0	2157	7	1	3	4864	4697	2028	
0	2158	7	1	3	4694	4866	2029	
0	2171	5	1	1	4825	
0	2172	6	1	2	4826	1919	
0	2173	5	1	1	4835	
0	2174	5	1	1	4830	
0	2175	5	1	1	4802	
0	2176	5	1	1	4840	
0	2177	7	1	3	4876	4707	2040	
0	2178	7	1	3	4704	4880	2041	
0	2194	5	2	1	4775	
0	2197	5	2	1	4893	
0	2200	5	1	1	4749	
0	2219	6	2	2	2031	2030	
0	2234	5	1	1	4811	
0	2235	5	1	1	4807	
0	2236	5	1	1	4820	
0	2237	5	1	1	4816	
0	2250	7	16	3	3943	4921	2119	
3	2266	3	0	2	1831	2126	
3	2269	3	0	2	2127	1832	
0	2291	3	2	2	2153	2154	
0	2294	3	2	2	2155	2156	
0	2297	4	1	2	2157	2032	
0	2298	4	1	2	2158	2033	
0	2300	5	1	1	4922	
0	2301	5	1	1	3899	
0	2302	6	1	2	3901	1519	
0	2303	5	1	1	3902	
0	2304	6	1	2	3905	1520	
0	2305	5	1	1	3906	
0	2306	6	1	2	3907	1521	
0	2307	5	1	1	3908	
0	2308	6	1	2	3920	1522	
0	2309	5	1	1	3921	
0	2310	6	1	2	3922	1523	
0	2311	5	1	1	3923	
0	2312	6	1	2	3991	1524	
0	2313	5	1	1	3992	
0	2314	6	1	2	3934	1525	
0	2315	5	1	1	3935	
0	2316	6	1	2	3936	1526	
0	2317	5	1	1	3937	
0	2318	6	1	2	4011	1527	
0	2319	5	1	1	4012	
0	2320	6	1	2	3940	1528	
0	2321	5	1	1	3941	
0	2322	6	1	2	4848	2171	
0	2323	6	1	2	4831	2173	
0	2324	6	1	2	4836	2174	
0	2325	6	1	2	4841	2175	
0	2326	6	1	2	4803	2176	
0	2327	4	1	2	2177	2042	
0	2328	4	1	2	2178	2043	
0	2329	6	1	2	4123	1572	
0	2330	5	1	1	4124	
0	2331	6	1	2	3948	1573	
0	2332	5	1	1	3949	
0	2333	6	1	2	3950	1574	
0	2334	5	1	1	3951	
0	2335	6	1	2	4231	1575	
0	2336	5	1	1	4232	
0	2337	6	1	2	4243	1576	
0	2338	5	1	1	4244	
0	2339	6	1	2	3954	1577	
0	2340	5	1	1	3955	
0	2354	6	1	2	4808	2234	
0	2355	6	1	2	4812	2235	
0	2356	6	1	2	4817	2236	
0	2357	6	1	2	4821	2237	
0	2358	7	1	2	4257	4294	
0	2359	5	28	1	3956	
0	2364	5	1	1	4898	
0	2365	5	1	1	4894	
0	2366	5	1	1	4904	
0	2367	5	1	1	3987	
0	2372	5	1	1	4899	
0	2373	5	1	1	4895	
0	2374	5	1	1	4905	
0	2375	5	1	1	4741	
0	2376	5	1	1	4906	
0	2377	5	4	1	3957	
0	2386	7	1	2	4258	4075	
0	2395	5	4	1	3958	
0	2400	6	1	2	3993	2300	
0	2403	5	1	1	4907	
0	2406	5	1	1	3994	
0	2407	6	1	2	4315	2303	
0	2408	6	1	2	4322	2305	
0	2409	6	1	2	4341	2307	
0	2410	6	1	2	4347	2309	
0	2411	6	1	2	4351	2311	
0	2412	6	1	2	4355	2313	
0	2413	6	1	2	4359	2315	
0	2414	6	1	2	4363	2317	
0	2415	6	1	2	4367	2319	
0	2416	6	1	2	4371	2321	
0	2417	6	3	2	2322	2172	
0	2421	6	3	2	2323	2324	
0	2425	6	4	2	2325	2326	
0	2428	6	1	2	4375	2330	
0	2429	6	1	2	4381	2332	
0	2430	6	1	2	4387	2334	
0	2431	6	1	2	4391	2336	
0	2432	6	1	2	4395	2338	
0	2433	6	1	2	4399	2340	
0	2452	5	1	1	3989	
0	2453	6	1	2	3990	2200	
0	2469	5	2	1	4259	
0	2484	6	2	2	2298	2297	
0	2487	6	2	2	2356	2357	
0	2490	6	2	2	2354	2355	
0	2493	6	2	2	2328	2327	
3	2496	3	0	2	2358	1814	
0	2503	6	1	2	4896	2364	
0	2504	6	1	2	4900	2365	
0	2510	6	1	2	4897	2372	
0	2511	6	1	2	4901	2373	
3	2521	3	0	2	1830	2386	
0	2528	6	1	2	4923	2406	
0	2531	5	2	1	4069	
0	2534	5	2	1	4077	
0	2544	6	1	2	2302	2407	
0	2545	6	1	2	2304	2408	
0	2546	6	1	2	2306	2409	
0	2547	6	1	2	2308	2410	
0	2548	6	1	2	2310	2411	
0	2549	6	1	2	2312	2412	
0	2550	6	1	2	2314	2413	
0	2551	6	1	2	2316	2414	
0	2552	6	1	2	2318	2415	
0	2553	6	1	2	2320	2416	
0	2563	6	1	2	2329	2428	
0	2564	6	1	2	2331	2429	
0	2565	6	1	2	2333	2430	
0	2566	6	1	2	2335	2431	
0	2567	6	1	2	2337	2432	
0	2568	6	1	2	2339	2433	
0	2579	6	1	2	4750	2452	
0	2607	7	1	2	4797	4217	
0	2608	7	1	2	4827	4218	
0	2609	7	1	2	4832	4219	
0	2610	7	1	2	4837	4220	
0	2611	7	1	2	4776	3959	
0	2612	7	1	2	4783	3960	
0	2613	6	3	2	2503	2504	
0	2617	5	1	1	4273	
0	2618	6	1	2	4274	2366	
0	2619	6	1	2	4285	2367	
0	2620	5	1	1	4286	
0	2621	5	2	1	4260	
0	2624	6	3	2	2510	2511	
0	2628	5	1	1	4275	
0	2629	6	1	2	4276	2374	
0	2630	5	1	1	4277	
0	2631	7	1	2	4777	3961	
0	2632	7	1	2	4784	3962	
0	2633	7	1	2	4798	4233	
0	2634	7	1	2	4828	4234	
0	2635	7	1	2	4833	4235	
0	2636	7	1	2	4838	4236	
0	2638	5	4	1	3963	
0	2645	5	1	1	4287	
0	2646	5	4	1	3964	
0	2652	6	1	2	2528	2400	
0	2655	5	1	1	4278	
0	2656	5	1	1	4288	
0	2663	5	1	1	4263	
0	2664	6	1	2	4264	2301	
0	2665	5	1	1	2553	
0	2666	5	1	1	2552	
0	2667	5	1	1	2551	
0	2668	5	1	1	2550	
0	2669	5	1	1	2549	
0	2670	5	1	1	2548	
0	2671	5	1	1	2547	
0	2672	5	1	1	2546	
0	2673	5	1	1	2545	
0	2674	5	1	1	2544	
0	2675	5	1	1	2568	
0	2676	5	1	1	2567	
0	2677	5	1	1	2566	
0	2678	5	1	1	2565	
0	2679	5	1	1	2564	
0	2680	5	1	1	2563	
0	2681	5	2	1	4245	
0	2684	5	2	1	4248	
0	2693	5	1	1	4269	
0	2694	6	1	2	4270	1807	
0	2695	5	1	1	3973	
0	2696	5	1	1	3969	
0	2697	5	1	1	3979	
0	2698	5	1	1	4305	
0	2699	5	1	1	3974	
0	2700	5	1	1	3970	
0	2701	5	1	1	3980	
0	2702	5	1	1	4306	
0	2703	6	2	2	2579	2453	
0	2706	5	1	1	4255	
0	2707	5	1	1	4265	
0	2708	5	1	1	4267	
0	2709	7	1	2	4078	4271	
0	2710	7	1	2	4070	4283	
0	2719	6	1	2	4908	2617	
0	2720	6	1	2	3988	2620	
0	2726	6	1	2	4909	2628	
0	2743	5	1	1	2652	
0	2747	6	1	2	3900	2663	
0	2748	7	1	5	2665	2666	2667	2668	2669	
0	2749	7	1	5	2670	2671	2672	2673	2674	
0	2750	7	1	2	2034	2675	
0	2751	7	1	5	2676	2677	2678	2679	2680	
0	2760	6	1	2	4727	2693	
0	2771	6	1	2	3971	2695	
0	2772	6	1	2	3975	2696	
0	2773	6	1	2	4307	2697	
0	2774	6	1	2	3981	2698	
0	2775	6	1	2	3972	2699	
0	2776	6	1	2	3976	2700	
0	2777	6	1	2	4308	2701	
0	2778	6	1	2	3982	2702	
0	2781	6	1	2	4268	2707	
0	2782	6	1	2	4266	2708	
0	2783	3	1	2	2709	4272	
0	2784	3	1	2	2710	4284	
0	2789	7	1	2	4778	4325	
0	2790	7	1	2	4785	4326	
0	2791	7	1	2	4789	4327	
0	2792	7	1	2	4793	4328	
0	2793	5	2	1	4309	
0	2796	6	3	2	2719	2618	
0	2800	6	4	2	2619	2720	
0	2803	5	2	1	4318	
0	2806	6	4	2	2726	2629	
0	2809	7	1	2	4779	4329	
0	2810	7	1	2	4786	4330	
0	2811	7	1	2	4790	4331	
0	2812	7	1	2	4794	4332	
3	2817	7	0	2	2743	14	
0	2826	6	2	2	2747	2664	
0	2829	7	1	2	2748	2749	
0	2830	7	1	2	2750	2751	
0	2837	5	1	1	4251	
0	2838	5	1	1	4252	
0	2839	7	1	3	4249	4246	4253	
0	2840	7	1	3	4335	4333	4254	
0	2841	6	2	2	2760	2694	
0	2874	6	2	2	2773	2774	
0	2877	6	2	2	2771	2772	
0	2880	5	1	1	4344	
0	2881	6	1	2	4345	2706	
0	2882	6	2	2	2777	2778	
0	2885	6	2	2	2775	2776	
0	2888	6	2	2	2781	2782	
3	2891	6	0	2	2783	2784	
0	2894	7	1	2	2607	3995	
0	2895	7	1	2	2608	3996	
0	2896	7	1	2	2609	3997	
0	2897	7	1	2	2610	3998	
0	2898	3	1	2	2789	2611	
0	2899	3	1	2	2790	2612	
0	2900	7	1	2	2791	3883	
0	2901	7	1	2	2792	3884	
0	2914	3	1	2	2809	2631	
0	2915	3	1	2	2810	2632	
0	2916	7	1	2	2811	3885	
0	2917	7	1	2	2812	3886	
0	2918	7	1	2	2633	3999	
0	2919	7	1	2	2634	4000	
0	2920	7	1	2	2635	4001	
0	2921	7	1	2	2636	4002	
3	2931	7	0	3	2829	2830	1302	
0	2938	7	1	3	4334	4250	2837	
0	2939	7	1	3	4247	4336	2838	
0	2963	6	1	2	4256	2880	
3	2970	5	0	1	4423	
3	2971	5	0	1	4421	
0	2972	5	3	1	2894	
0	2975	5	3	1	2895	
0	2978	5	3	1	2896	
0	2981	5	3	1	2897	
0	2984	7	1	2	2898	3887	
0	2985	7	1	2	2899	3888	
0	2986	5	3	1	2900	
0	2989	5	3	1	2901	
0	2992	5	2	1	4408	
0	3007	7	1	2	4316	4133	
0	3008	7	1	2	2914	3889	
0	3009	7	1	2	2915	3890	
0	3010	5	3	1	2916	
0	3013	5	3	1	2917	
0	3016	5	3	1	2918	
0	3019	5	3	1	2919	
0	3022	5	3	1	2920	
0	3025	5	3	1	2921	
0	3028	5	1	1	2817	
0	3029	7	1	2	4317	4134	
0	3030	5	4	1	4135	
0	3035	7	1	2	4323	4136	
0	3036	7	1	2	4342	4137	
0	3037	7	1	2	4348	4138	
0	3039	5	4	1	4139	
0	3044	7	1	2	4324	4140	
0	3045	7	1	2	4343	4141	
0	3046	7	1	2	4349	4142	
0	3047	4	1	2	2938	2839	
0	3048	4	1	2	2939	2840	
0	3049	5	1	1	4435	
0	3050	5	2	1	4143	
0	3053	7	1	2	4352	4144	
0	3054	7	1	2	4356	4145	
0	3055	7	1	2	4360	4146	
0	3056	7	1	2	4364	4147	
0	3057	7	1	2	4368	4148	
0	3058	7	1	2	4372	4149	
0	3059	7	1	2	4376	4150	
0	3060	7	1	2	4382	4151	
0	3061	5	2	1	4152	
0	3064	7	1	2	4353	4153	
0	3065	7	1	2	4357	4154	
0	3066	7	1	2	4361	4155	
0	3067	7	1	2	4365	4156	
0	3068	7	1	2	4369	4157	
0	3069	7	1	2	4373	4158	
0	3070	7	1	2	4377	4159	
0	3071	7	1	2	4383	4160	
0	3072	5	1	1	4427	
0	3073	5	1	1	4429	
0	3074	5	1	1	4431	
0	3075	5	1	1	4433	
0	3076	6	2	2	2881	2963	
3	3079	5	0	1	2931	
0	3088	5	3	1	2984	
0	3091	5	3	1	2985	
0	3110	5	3	1	3008	
0	3113	5	3	1	3009	
0	3137	7	3	2	3055	3891	
0	3140	7	3	2	3056	3892	
0	3143	7	3	2	3057	4003	
0	3146	7	3	2	3058	4004	
0	3149	7	3	2	3059	4005	
0	3152	7	3	2	3060	4006	
0	3157	7	3	2	3066	3893	
0	3160	7	3	2	3067	3894	
0	3163	7	3	2	3068	4007	
0	3166	7	3	2	3069	4008	
0	3169	7	3	2	3070	4009	
0	3172	7	3	2	3071	4010	
0	3175	6	1	2	4430	3072	
0	3176	6	1	2	4428	3073	
0	3177	6	1	2	4434	3074	
0	3178	6	1	2	4432	3075	
0	3180	6	2	2	3048	3047	
0	3187	5	1	1	4411	
0	3188	5	1	1	4412	
0	3189	5	1	1	4417	
0	3190	5	1	1	4418	
0	3191	7	1	3	4409	4310	4413	
0	3192	7	1	3	4455	4406	4414	
0	3193	7	1	3	4319	4261	4419	
0	3194	7	1	3	4415	4312	4420	
0	3195	6	1	2	4489	2375	
0	3196	5	1	1	4490	
0	3197	7	1	2	4378	4475	
0	3208	7	1	2	4379	4481	
0	3215	7	1	2	4384	4476	
0	3216	7	1	2	4388	4477	
0	3217	7	1	2	4392	4478	
0	3218	7	1	2	4385	4482	
0	3219	7	1	2	4389	4483	
0	3220	7	1	2	4393	4484	
0	3222	7	1	2	4396	4485	
0	3223	7	1	2	4400	4486	
0	3230	7	1	2	4397	4487	
0	3231	7	1	2	4401	4488	
0	3238	6	2	2	3175	3176	
0	3241	6	2	2	3177	3178	
0	3281	7	1	3	4407	4410	3187	
0	3282	7	1	3	4311	4456	3188	
0	3283	7	1	3	4313	4320	3189	
0	3284	7	1	3	4262	4416	3190	
0	3286	6	1	2	4742	3196	
0	3288	3	1	2	3197	3007	
0	3289	6	1	2	4607	3049	
0	3291	7	1	2	4570	4446	
0	3293	7	1	2	4567	4443	
0	3295	7	1	2	4564	4440	
0	3296	7	1	2	4437	4551	
0	3299	7	1	2	4548	4452	
0	3301	7	1	2	4545	4449	
0	3302	3	1	2	3208	3029	
0	3304	7	1	2	4601	4472	
0	3306	7	1	2	4595	4469	
0	3308	7	1	2	4592	4466	
0	3309	7	1	2	4463	4589	
0	3312	7	1	2	4576	4460	
0	3314	7	1	2	4573	4457	
0	3315	3	3	2	3215	3035	
0	3318	3	3	2	3216	3036	
0	3321	3	3	2	3217	3037	
0	3324	3	3	2	3218	3044	
0	3327	3	3	2	3219	3045	
0	3330	3	3	2	3220	3046	
0	3333	5	1	1	4608	
0	3334	3	1	2	3222	3053	
0	3335	3	1	2	3223	3054	
0	3336	3	1	2	3230	3064	
0	3337	3	1	2	3231	3065	
0	3400	6	1	2	3195	3286	
0	3401	4	1	2	3281	3191	
0	3402	4	1	2	3282	3192	
0	3403	4	1	2	3283	3193	
0	3404	4	1	2	3284	3194	
0	3405	5	1	1	4642	
0	3406	5	1	1	4644	
0	3409	7	1	2	3288	4902	
0	3410	6	1	2	4436	3333	
0	3412	5	1	1	4447	
0	3414	5	1	1	4444	
0	3416	5	1	1	4441	
0	3418	5	1	1	4438	
0	3420	5	1	1	4453	
0	3422	5	1	1	4450	
0	3428	7	1	2	3302	4903	
0	3430	5	1	1	4473	
0	3432	5	1	1	4470	
0	3434	5	1	1	4467	
0	3436	5	1	1	4464	
0	3438	5	1	1	4461	
0	3440	5	1	1	4458	
0	3450	7	3	2	3334	3895	
0	3453	7	3	2	3335	3896	
0	3456	7	3	2	3336	3897	
0	3459	7	3	2	3337	3898	
0	3478	7	1	2	3400	4295	
0	3479	7	1	2	4659	4279	
0	3480	7	1	2	4656	4910	
0	3481	6	1	2	3410	3289	
0	3482	5	1	1	4571	
0	3483	6	1	2	4572	3412	
0	3484	5	1	1	4568	
0	3485	6	1	2	4569	3414	
0	3486	5	1	1	4565	
0	3487	6	1	2	4566	3416	
0	3488	5	1	1	4552	
0	3489	6	1	2	4553	3418	
0	3490	5	1	1	4549	
0	3491	6	1	2	4550	3420	
0	3492	5	1	1	4546	
0	3493	6	1	2	4547	3422	
0	3494	5	1	1	4504	
0	3496	5	1	1	4491	
0	3498	7	1	2	4662	4289	
0	3499	7	1	2	4668	4280	
0	3500	7	1	2	4665	4911	
0	3501	5	1	1	4602	
0	3502	6	1	2	4603	3430	
0	3503	5	1	1	4596	
0	3504	6	1	2	4597	3432	
0	3505	5	1	1	4593	
0	3506	6	1	2	4594	3434	
0	3507	5	1	1	4590	
0	3508	6	1	2	4591	3436	
0	3509	5	1	1	4577	
0	3510	6	1	2	4578	3438	
0	3511	5	1	1	4574	
0	3512	6	1	2	4575	3440	
0	3513	5	1	1	4522	
0	3515	5	1	1	4519	
0	3517	7	1	2	4671	4290	
0	3522	6	2	2	3402	3401	
0	3525	6	2	2	3404	3403	
3	3546	3	0	2	3478	1813	
0	3551	5	1	1	3481	
0	3552	6	1	2	4448	3482	
0	3553	6	1	2	4445	3484	
0	3554	6	1	2	4442	3486	
0	3555	6	1	2	4439	3488	
0	3556	6	1	2	4454	3490	
0	3557	6	1	2	4451	3492	
0	3558	7	1	2	4679	4505	
0	3559	7	1	2	4676	4492	
0	3563	6	1	2	4474	3501	
0	3564	6	1	2	4471	3503	
0	3565	6	1	2	4468	3505	
0	3566	6	1	2	4465	3507	
0	3567	6	1	2	4462	3509	
0	3568	6	1	2	4459	3511	
0	3569	7	1	2	4685	4523	
0	3570	7	1	2	4682	4520	
0	3592	5	1	1	4674	
0	3593	6	1	2	4675	3405	
0	3594	5	1	1	4517	
0	3595	6	1	2	4518	3406	
0	3596	5	1	1	4660	
0	3597	6	1	2	4661	2630	
0	3598	6	1	2	4657	2376	
0	3599	5	1	1	4658	
3	3600	7	0	2	3551	4425	
0	3603	6	4	2	3552	3483	
0	3608	6	3	2	3553	3485	
0	3612	6	2	2	3554	3487	
0	3615	6	1	2	3555	3489	
0	3616	6	5	2	3556	3491	
0	3622	6	4	2	3557	3493	
0	3629	5	1	1	4663	
0	3630	6	1	2	4664	2645	
0	3631	5	1	1	4669	
0	3632	6	1	2	4670	2655	
0	3633	6	1	2	4666	2403	
0	3634	5	1	1	4667	
0	3635	6	4	2	3563	3502	
0	3640	6	3	2	3564	3504	
0	3644	6	2	2	3565	3506	
0	3647	6	1	2	3566	3508	
0	3648	6	5	2	3567	3510	
0	3654	6	4	2	3568	3512	
0	3661	5	1	1	4672	
0	3662	6	1	2	4673	2656	
0	3667	6	1	2	4643	3592	
0	3668	6	1	2	4645	3594	
0	3669	6	1	2	4281	3596	
0	3670	6	1	2	4912	3599	
0	3691	5	1	1	4680	
0	3692	6	1	2	4681	3494	
0	3693	5	1	1	4677	
0	3694	6	1	2	4678	3496	
0	3695	6	1	2	4291	3629	
0	3696	6	1	2	4282	3631	
0	3697	6	1	2	4913	3634	
0	3716	5	1	1	4686	
0	3717	6	1	2	4687	3513	
0	3718	5	1	1	4683	
0	3719	6	1	2	4684	3515	
0	3720	6	1	2	4292	3661	
0	3721	6	1	2	3667	3593	
0	3722	6	1	2	3668	3595	
0	3723	6	2	2	3669	3597	
0	3726	6	1	2	3670	3598	
0	3727	5	1	1	3600	
0	3728	6	1	2	4506	3691	
0	3729	6	1	2	4493	3693	
0	3730	6	1	2	3695	3630	
0	3731	7	1	4	4860	3615	4871	4712	
0	3732	7	1	2	4713	3293	
0	3733	7	1	3	4861	4714	3295	
0	3734	7	1	4	4872	4715	3296	4862	
0	3735	7	1	2	4883	3301	
0	3736	7	1	3	4720	4884	3558	
0	3737	6	2	2	3696	3632	
0	3740	6	1	2	3697	3633	
0	3741	6	1	2	4524	3716	
0	3742	6	1	2	4521	3718	
0	3743	6	1	2	3720	3662	
0	3744	7	1	4	4735	3647	4743	4731	
0	3745	7	1	2	4732	3306	
0	3746	7	1	3	4736	4733	3308	
0	3747	7	1	4	4744	4734	3309	4737	
0	3748	7	1	2	4751	3314	
0	3749	7	1	3	4761	4752	3569	
0	3750	5	1	1	3721	
0	3753	7	1	2	3722	4076	
0	3754	6	3	2	3728	3692	
0	3758	6	2	2	3729	3694	
0	3761	5	1	1	3731	
0	3762	3	2	4	3291	3732	3733	3734	
0	3767	6	3	2	3741	3717	
0	3771	6	2	2	3742	3719	
0	3774	5	1	1	3744	
0	3775	3	2	4	3304	3745	3746	3747	
0	3778	7	1	2	4822	3480	
0	3779	7	1	3	3726	4823	3409	
3	3780	3	0	2	2125	3753	
3	3790	7	0	2	3750	4426	
0	3793	7	1	2	4842	3500	
0	3794	7	1	3	3740	4843	3428	
0	3802	3	1	3	3479	3778	3779	
0	3805	5	1	1	4851	
0	3806	7	1	5	4721	3730	4844	4885	4849	
0	3807	7	1	4	4845	4886	3559	4722	
0	3808	7	1	5	4850	4846	4887	3498	4723	
0	3811	3	1	3	3499	3793	3794	
0	3812	5	1	1	4858	
0	3813	7	1	5	4762	3743	4853	4753	4856	
0	3814	7	1	4	4854	4754	3570	4763	
0	3815	7	1	5	4857	4855	4755	3517	4764	
0	3816	3	1	5	3299	3735	3736	3807	3808	
0	3817	7	1	2	3806	3802	
0	3818	6	1	2	3805	3761	
0	3819	5	1	1	3790	
0	3820	3	1	5	3312	3748	3749	3814	3815	
0	3821	7	1	2	3813	3811	
0	3822	6	1	2	3812	3774	
0	3823	3	2	2	3816	3817	
0	3826	7	1	3	3727	3819	4424	
0	3827	3	2	2	3820	3821	
0	3834	5	1	1	4867	
0	3835	7	1	2	3818	4868	
0	3836	5	1	1	4869	
0	3837	7	1	2	3822	4870	
0	3838	7	1	2	4852	3834	
0	3839	7	1	2	4859	3836	
0	3840	3	2	2	3838	3835	
3	3843	3	0	2	3839	3837	
0	3852	6	2	2	4877	4873	
0	3857	7	1	2	4878	4881	
0	3858	7	1	2	4882	4874	
0	3859	3	2	2	3857	3858	
0	3864	5	2	1	4479	
0	3869	7	1	2	4480	4888	
0	3870	3	2	2	3869	4889	
3	3875	5	0	1	4890	
0	3876	7	1	3	4422	3028	4891	
3	3877	7	0	3	3826	3876	4730	
3	3882	5	0	1	3877	
2	3883	1	8			
2	3884	1	8			
2	3885	1	8			
2	3886	1	8			
2	3887	1	8			
2	3888	1	8			
2	3889	1	8			
2	3890	1	8			
2	3891	1	8			
2	3892	1	8			
2	3893	1	8			
2	3894	1	8			
2	3895	1	8			
2	3896	1	8			
2	3897	1	8			
2	3898	1	8			
2	3899	1	2049			
2	3900	1	2049			
2	3901	1	2052			
2	3902	1	2052			
2	3903	1	11			
2	3904	1	11			
2	3905	1	2055			
2	3906	1	2055			
2	3907	1	2058			
2	3908	1	2058			
2	3909	1	16			
2	3910	1	16			
2	3911	1	16			
2	3912	1	16			
2	3913	1	16			
2	3914	1	16			
2	3915	1	16			
2	3916	1	16			
2	3917	1	16			
2	3918	1	16			
2	3919	1	16			
2	3920	1	2061			
2	3921	1	2061			
2	3922	1	2064			
2	3923	1	2064			
2	3924	1	29			
2	3925	1	29			
2	3926	1	29			
2	3927	1	29			
2	3928	1	29			
2	3929	1	29			
2	3930	1	29			
2	3931	1	29			
2	3932	1	29			
2	3933	1	29			
2	3934	1	2070			
2	3935	1	2070			
2	3936	1	2073			
2	3937	1	2073			
2	3938	1	37			
2	3939	1	37			
2	3940	1	2079			
2	3941	1	2079			
2	3942	1	40			
2	3943	1	40			
2	3944	1	44			
2	3945	1	44			
2	3946	1	57			
2	3947	1	57			
2	3948	1	2098			
2	3949	1	2098			
2	3950	1	2101			
2	3951	1	2101			
2	3952	1	69			
2	3953	1	69			
2	3954	1	2110			
2	3955	1	2110			
2	3956	1	2113			
2	3957	1	2113			
2	3958	1	2113			
2	3959	1	2113			
2	3960	1	2113			
2	3961	1	2113			
2	3962	1	2113			
2	3963	1	2113			
2	3964	1	2113			
2	3965	1	82			
2	3966	1	82			
2	3967	1	96			
2	3968	1	96			
2	3969	1	2141			
2	3970	1	2141			
2	3971	1	2141			
2	3972	1	2141			
2	3973	1	2144			
2	3974	1	2144			
2	3975	1	2144			
2	3976	1	2144			
2	3977	1	108			
2	3978	1	108			
2	3979	1	2150			
2	3980	1	2150			
2	3981	1	2150			
2	3982	1	2150			
2	3983	1	120			
2	3984	1	120			
2	3985	1	132			
2	3986	1	132			
2	3987	1	2194			
2	3988	1	2194			
2	3989	1	2197			
2	3990	1	2197			
2	3991	1	2067			
2	3992	1	2067			
2	3993	1	2219			
2	3994	1	2219			
2	3995	1	2250			
2	3996	1	2250			
2	3997	1	2250			
2	3998	1	2250			
2	3999	1	2250			
2	4000	1	2250			
2	4001	1	2250			
2	4002	1	2250			
2	4003	1	2250			
2	4004	1	2250			
2	4005	1	2250			
2	4006	1	2250			
2	4007	1	2250			
2	4008	1	2250			
2	4009	1	2250			
2	4010	1	2250			
2	4011	1	2076			
2	4012	1	2076			
2	4013	1	224			
2	4014	1	224			
2	4015	1	227			
2	4016	1	227			
2	4017	1	227			
2	4018	1	227			
2	4019	1	227			
2	4020	1	227			
2	4021	1	227			
2	4022	1	227			
2	4023	1	227			
2	4024	1	227			
2	4025	1	227			
2	4026	1	227			
2	4027	1	227			
2	4028	1	227			
2	4029	1	227			
2	4030	1	227			
2	4031	1	227			
2	4032	1	227			
2	4033	1	227			
2	4034	1	227			
2	4035	1	227			
2	4036	1	227			
2	4037	1	231			
2	4038	1	231			
2	4039	1	234			
2	4040	1	234			
2	4041	1	234			
2	4042	1	234			
2	4043	1	234			
2	4044	1	234			
2	4045	1	234			
2	4046	1	234			
2	4047	1	234			
2	4048	1	234			
2	4049	1	234			
2	4050	1	234			
2	4051	1	234			
2	4052	1	234			
2	4053	1	234			
2	4054	1	234			
2	4055	1	234			
2	4056	1	234			
2	4057	1	234			
2	4058	1	234			
2	4059	1	234			
2	4060	1	234			
2	4061	1	237			
2	4062	1	237			
2	4063	1	237			
2	4064	1	237			
2	4065	1	241			
2	4066	1	241			
2	4067	1	241			
2	4068	1	241			
2	4069	1	2291			
2	4070	1	2291			
2	4071	1	246			
2	4072	1	246			
2	4073	1	246			
2	4074	1	246			
2	4075	1	246			
2	4076	1	246			
2	4077	1	2294			
2	4078	1	2294			
2	4079	1	256			
2	4080	1	256			
2	4081	1	256			
2	4082	1	259			
2	4083	1	259			
2	4084	1	259			
2	4085	1	263			
2	4086	1	263			
2	4087	1	263			
2	4088	1	266			
2	4089	1	266			
2	4090	1	266			
2	4091	1	269			
2	4092	1	269			
2	4093	1	269			
2	4094	1	272			
2	4095	1	272			
2	4096	1	272			
2	4097	1	275			
2	4098	1	275			
2	4099	1	275			
2	4100	1	278			
2	4101	1	278			
2	4102	1	278			
2	4103	1	281			
2	4104	1	281			
2	4105	1	281			
2	4106	1	284			
2	4107	1	284			
2	4108	1	284			
2	4109	1	287			
2	4110	1	287			
2	4111	1	287			
2	4112	1	294			
2	4113	1	294			
2	4114	1	294			
2	4115	1	297			
2	4116	1	297			
2	4117	1	297			
2	4118	1	297			
2	4119	1	301			
2	4120	1	301			
2	4121	1	301			
2	4122	1	301			
2	4123	1	2095			
2	4124	1	2095			
2	4125	1	305			
2	4126	1	305			
2	4127	1	305			
2	4128	1	305			
2	4129	1	309			
2	4130	1	309			
2	4131	1	309			
2	4132	1	309			
2	4133	1	2359			
2	4134	1	2359			
2	4135	1	2359			
2	4136	1	2359			
2	4137	1	2359			
2	4138	1	2359			
2	4139	1	2359			
2	4140	1	2359			
2	4141	1	2359			
2	4142	1	2359			
2	4143	1	2359			
2	4144	1	2359			
2	4145	1	2359			
2	4146	1	2359			
2	4147	1	2359			
2	4148	1	2359			
2	4149	1	2359			
2	4150	1	2359			
2	4151	1	2359			
2	4152	1	2359			
2	4153	1	2359			
2	4154	1	2359			
2	4155	1	2359			
2	4156	1	2359			
2	4157	1	2359			
2	4158	1	2359			
2	4159	1	2359			
2	4160	1	2359			
2	4161	1	313			
2	4162	1	313			
2	4163	1	313			
2	4164	1	316			
2	4165	1	316			
2	4166	1	316			
2	4167	1	319			
2	4168	1	319			
2	4169	1	319			
2	4170	1	319			
2	4171	1	319			
2	4172	1	319			
2	4173	1	319			
2	4174	1	319			
2	4175	1	319			
2	4176	1	319			
2	4177	1	319			
2	4178	1	319			
2	4179	1	319			
2	4180	1	319			
2	4181	1	319			
2	4182	1	319			
2	4183	1	319			
2	4184	1	319			
2	4185	1	319			
2	4186	1	319			
2	4187	1	319			
2	4188	1	319			
2	4189	1	322			
2	4190	1	322			
2	4191	1	322			
2	4192	1	322			
2	4193	1	322			
2	4194	1	322			
2	4195	1	322			
2	4196	1	322			
2	4197	1	322			
2	4198	1	322			
2	4199	1	322			
2	4200	1	322			
2	4201	1	322			
2	4202	1	322			
2	4203	1	322			
2	4204	1	322			
2	4205	1	322			
2	4206	1	322			
2	4207	1	322			
2	4208	1	322			
2	4209	1	322			
2	4210	1	322			
2	4211	1	325			
2	4212	1	325			
2	4213	1	328			
2	4214	1	328			
2	4215	1	331			
2	4216	1	331			
2	4217	1	2377			
2	4218	1	2377			
2	4219	1	2377			
2	4220	1	2377			
2	4221	1	334			
2	4222	1	334			
2	4223	1	337			
2	4224	1	337			
2	4225	1	340			
2	4226	1	340			
2	4227	1	343			
2	4228	1	343			
2	4229	1	346			
2	4230	1	346			
2	4231	1	2104			
2	4232	1	2104			
2	4233	1	2395			
2	4234	1	2395			
2	4235	1	2395			
2	4236	1	2395			
2	4237	1	349			
2	4238	1	349			
2	4239	1	352			
2	4240	1	352			
2	4241	1	355			
2	4242	1	355			
2	4243	1	2107			
2	4244	1	2107			
2	4245	1	2417			
2	4246	1	2417			
2	4247	1	2417			
2	4248	1	2421			
2	4249	1	2421			
2	4250	1	2421			
2	4251	1	2425			
2	4252	1	2425			
2	4253	1	2425			
2	4254	1	2425			
2	4255	1	2469			
2	4256	1	2469			
2	4257	1	2120			
2	4258	1	2120			
2	4259	1	2120			
2	4260	1	2120			
2	4261	1	2120			
2	4262	1	2120			
2	4263	1	2484			
2	4264	1	2484			
2	4265	1	2487			
2	4266	1	2487			
2	4267	1	2490			
2	4268	1	2490			
2	4269	1	2493			
2	4270	1	2493			
2	4271	1	2534			
2	4272	1	2534			
2	4273	1	2128			
2	4274	1	2128			
2	4275	1	2128			
2	4276	1	2128			
2	4277	1	2128			
2	4278	1	2128			
2	4279	1	2128			
2	4280	1	2128			
2	4281	1	2128			
2	4282	1	2128			
2	4283	1	2531			
2	4284	1	2531			
2	4285	1	2135			
2	4286	1	2135			
2	4287	1	2135			
2	4288	1	2135			
2	4289	1	2135			
2	4290	1	2135			
2	4291	1	2135			
2	4292	1	2135			
2	4293	1	533			
2	4294	1	533			
2	4295	1	533			
2	4296	1	537			
2	4297	1	537			
2	4298	1	537			
2	4299	1	537			
2	4300	1	537			
2	4301	1	544			
2	4302	1	544			
2	4303	1	547			
2	4304	1	547			
2	4305	1	2147			
2	4306	1	2147			
2	4307	1	2147			
2	4308	1	2147			
2	4309	1	2613			
2	4310	1	2613			
2	4311	1	2613			
2	4312	1	2621			
2	4313	1	2621			
2	4314	1	574			
2	4315	1	574			
2	4316	1	574			
2	4317	1	574			
2	4318	1	2624			
2	4319	1	2624			
2	4320	1	2624			
2	4321	1	578			
2	4322	1	578			
2	4323	1	578			
2	4324	1	578			
2	4325	1	2638			
2	4326	1	2638			
2	4327	1	2638			
2	4328	1	2638			
2	4329	1	2646			
2	4330	1	2646			
2	4331	1	2646			
2	4332	1	2646			
2	4333	1	2681			
2	4334	1	2681			
2	4335	1	2684			
2	4336	1	2684			
2	4337	1	651			
2	4338	1	651			
2	4339	1	651			
2	4340	1	655			
2	4341	1	655			
2	4342	1	655			
2	4343	1	655			
2	4344	1	2703			
2	4345	1	2703			
2	4346	1	659			
2	4347	1	659			
2	4348	1	659			
2	4349	1	659			
2	4350	1	663			
2	4351	1	663			
2	4352	1	663			
2	4353	1	663			
2	4354	1	667			
2	4355	1	667			
2	4356	1	667			
2	4357	1	667			
2	4358	1	671			
2	4359	1	671			
2	4360	1	671			
2	4361	1	671			
2	4362	1	675			
2	4363	1	675			
2	4364	1	675			
2	4365	1	675			
2	4366	1	679			
2	4367	1	679			
2	4368	1	679			
2	4369	1	679			
2	4370	1	683			
2	4371	1	683			
2	4372	1	683			
2	4373	1	683			
2	4374	1	687			
2	4375	1	687			
2	4376	1	687			
2	4377	1	687			
2	4378	1	687			
2	4379	1	687			
2	4380	1	705			
2	4381	1	705			
2	4382	1	705			
2	4383	1	705			
2	4384	1	705			
2	4385	1	705			
2	4386	1	711			
2	4387	1	711			
2	4388	1	711			
2	4389	1	711			
2	4390	1	715			
2	4391	1	715			
2	4392	1	715			
2	4393	1	715			
2	4394	1	719			
2	4395	1	719			
2	4396	1	719			
2	4397	1	719			
2	4398	1	723			
2	4399	1	723			
2	4400	1	723			
2	4401	1	723			
2	4402	1	727			
2	4403	1	727			
2	4404	1	730			
2	4405	1	730			
2	4406	1	2793			
2	4407	1	2793			
2	4408	1	2796			
2	4409	1	2796			
2	4410	1	2796			
2	4411	1	2800			
2	4412	1	2800			
2	4413	1	2800			
2	4414	1	2800			
2	4415	1	2803			
2	4416	1	2803			
2	4417	1	2806			
2	4418	1	2806			
2	4419	1	2806			
2	4420	1	2806			
2	4421	1	2826			
2	4422	1	2826			
2	4423	1	2841			
2	4424	1	2841			
2	4425	1	800			
2	4426	1	800			
2	4427	1	2874			
2	4428	1	2874			
2	4429	1	2877			
2	4430	1	2877			
2	4431	1	2882			
2	4432	1	2882			
2	4433	1	2885			
2	4434	1	2885			
2	4435	1	2888			
2	4436	1	2888			
2	4437	1	2972			
2	4438	1	2972			
2	4439	1	2972			
2	4440	1	2975			
2	4441	1	2975			
2	4442	1	2975			
2	4443	1	2978			
2	4444	1	2978			
2	4445	1	2978			
2	4446	1	2981			
2	4447	1	2981			
2	4448	1	2981			
2	4449	1	2986			
2	4450	1	2986			
2	4451	1	2986			
2	4452	1	2989			
2	4453	1	2989			
2	4454	1	2989			
2	4455	1	2992			
2	4456	1	2992			
2	4457	1	3010			
2	4458	1	3010			
2	4459	1	3010			
2	4460	1	3013			
2	4461	1	3013			
2	4462	1	3013			
2	4463	1	3016			
2	4464	1	3016			
2	4465	1	3016			
2	4466	1	3019			
2	4467	1	3019			
2	4468	1	3019			
2	4469	1	3022			
2	4470	1	3022			
2	4471	1	3022			
2	4472	1	3025			
2	4473	1	3025			
2	4474	1	3025			
2	4475	1	3030			
2	4476	1	3030			
2	4477	1	3030			
2	4478	1	3030			
2	4479	1	3859			
2	4480	1	3859			
2	4481	1	3039			
2	4482	1	3039			
2	4483	1	3039			
2	4484	1	3039			
2	4485	1	3050			
2	4486	1	3050			
2	4487	1	3061			
2	4488	1	3061			
2	4489	1	3076			
2	4490	1	3076			
2	4491	1	3088			
2	4492	1	3088			
2	4493	1	3088			
2	4494	1	1042			
2	4495	1	1042			
2	4496	1	1042			
2	4497	1	1042			
2	4498	1	1042			
2	4499	1	1042			
2	4500	1	1042			
2	4501	1	1042			
2	4502	1	1042			
2	4503	1	1042			
2	4504	1	3091			
2	4505	1	3091			
2	4506	1	3091			
2	4507	1	1053			
2	4508	1	1053			
2	4509	1	1053			
2	4510	1	1053			
2	4511	1	1053			
2	4512	1	1053			
2	4513	1	1053			
2	4514	1	1053			
2	4515	1	1053			
2	4516	1	1053			
2	4517	1	3525			
2	4518	1	3525			
2	4519	1	3110			
2	4520	1	3110			
2	4521	1	3110			
2	4522	1	3113			
2	4523	1	3113			
2	4524	1	3113			
2	4525	1	1075			
2	4526	1	1075			
2	4527	1	1075			
2	4528	1	1075			
2	4529	1	1075			
2	4530	1	1075			
2	4531	1	1075			
2	4532	1	1075			
2	4533	1	1075			
2	4534	1	1075			
2	4535	1	1086			
2	4536	1	1086			
2	4537	1	1086			
2	4538	1	1086			
2	4539	1	1086			
2	4540	1	1086			
2	4541	1	1086			
2	4542	1	1086			
2	4543	1	1086			
2	4544	1	1086			
2	4545	1	3137			
2	4546	1	3137			
2	4547	1	3137			
2	4548	1	3140			
2	4549	1	3140			
2	4550	1	3140			
2	4551	1	3143			
2	4552	1	3143			
2	4553	1	3143			
2	4554	1	1102			
2	4555	1	1102			
2	4556	1	1102			
2	4557	1	1102			
2	4558	1	1102			
2	4559	1	1102			
2	4560	1	1102			
2	4561	1	1102			
2	4562	1	1102			
2	4563	1	1102			
2	4564	1	3146			
2	4565	1	3146			
2	4566	1	3146			
2	4567	1	3149			
2	4568	1	3149			
2	4569	1	3149			
2	4570	1	3152			
2	4571	1	3152			
2	4572	1	3152			
2	4573	1	3157			
2	4574	1	3157			
2	4575	1	3157			
2	4576	1	3160			
2	4577	1	3160			
2	4578	1	3160			
2	4579	1	1113			
2	4580	1	1113			
2	4581	1	1113			
2	4582	1	1113			
2	4583	1	1113			
2	4584	1	1113			
2	4585	1	1113			
2	4586	1	1113			
2	4587	1	1113			
2	4588	1	1113			
2	4589	1	3163			
2	4590	1	3163			
2	4591	1	3163			
2	4592	1	3166			
2	4593	1	3166			
2	4594	1	3166			
2	4595	1	3169			
2	4596	1	3169			
2	4597	1	3169			
2	4598	1	1129			
2	4599	1	1129			
2	4600	1	1129			
2	4601	1	3172			
2	4602	1	3172			
2	4603	1	3172			
2	4604	1	1133			
2	4605	1	1133			
2	4606	1	1133			
2	4607	1	3180			
2	4608	1	3180			
2	4609	1	1137			
2	4610	1	1137			
2	4611	1	1137			
2	4612	1	1137			
2	4613	1	1146			
2	4614	1	1146			
2	4615	1	1146			
2	4616	1	1146			
2	4617	1	1146			
2	4618	1	1146			
2	4619	1	1146			
2	4620	1	1146			
2	4621	1	1146			
2	4622	1	1146			
2	4623	1	1157			
2	4624	1	1157			
2	4625	1	1157			
2	4626	1	1157			
2	4627	1	1157			
2	4628	1	1157			
2	4629	1	1157			
2	4630	1	1157			
2	4631	1	1157			
2	4632	1	1157			
2	4633	1	1173			
2	4634	1	1173			
2	4635	1	1173			
2	4636	1	1173			
2	4637	1	1178			
2	4638	1	1178			
2	4639	1	1178			
2	4640	1	1178			
2	4641	1	1178			
2	4642	1	3238			
2	4643	1	3238			
2	4644	1	3241			
2	4645	1	3241			
2	4646	1	1200			
2	4647	1	1200			
2	4648	1	1200			
2	4649	1	1200			
2	4650	1	1205			
2	4651	1	1205			
2	4652	1	1205			
2	4653	1	1205			
2	4654	1	1216			
2	4655	1	1216			
2	4656	1	3315			
2	4657	1	3315			
2	4658	1	3315			
2	4659	1	3318			
2	4660	1	3318			
2	4661	1	3318			
2	4662	1	3321			
2	4663	1	3321			
2	4664	1	3321			
2	4665	1	3324			
2	4666	1	3324			
2	4667	1	3324			
2	4668	1	3327			
2	4669	1	3327			
2	4670	1	3327			
2	4671	1	3330			
2	4672	1	3330			
2	4673	1	3330			
2	4674	1	3522			
2	4675	1	3522			
2	4676	1	3450			
2	4677	1	3450			
2	4678	1	3450			
2	4679	1	3453			
2	4680	1	3453			
2	4681	1	3453			
2	4682	1	3456			
2	4683	1	3456			
2	4684	1	3456			
2	4685	1	3459			
2	4686	1	3459			
2	4687	1	3459			
2	4688	1	1496			
2	4689	1	1496			
2	4690	1	1499			
2	4691	1	1499			
2	4692	1	1502			
2	4693	1	1502			
2	4694	1	1502			
2	4695	1	1506			
2	4696	1	1506			
2	4697	1	1506			
2	4698	1	1510			
2	4699	1	1510			
2	4700	1	1510			
2	4701	1	1510			
2	4702	1	1553			
2	4703	1	1553			
2	4704	1	1553			
2	4705	1	1557			
2	4706	1	1557			
2	4707	1	1557			
2	4708	1	1561			
2	4709	1	1561			
2	4710	1	1561			
2	4711	1	1561			
2	4712	1	3603			
2	4713	1	3603			
2	4714	1	3603			
2	4715	1	3603			
2	4716	1	1578			
2	4717	1	1578			
2	4718	1	1582			
2	4719	1	1582			
2	4720	1	3622			
2	4721	1	3622			
2	4722	1	3622			
2	4723	1	3622			
2	4724	1	1585			
2	4725	1	1585			
2	4726	1	1588			
2	4727	1	1588			
2	4728	1	1591			
2	4729	1	1591			
2	4730	1	1591			
2	4731	1	3635			
2	4732	1	3635			
2	4733	1	3635			
2	4734	1	3635			
2	4735	1	3640			
2	4736	1	3640			
2	4737	1	3640			
2	4738	1	1596			
2	4739	1	1596			
2	4740	1	1596			
2	4741	1	1596			
2	4742	1	1596			
2	4743	1	3644			
2	4744	1	3644			
2	4745	1	1600			
2	4746	1	1600			
2	4747	1	1600			
2	4748	1	1600			
2	4749	1	1600			
2	4750	1	1600			
2	4751	1	3648			
2	4752	1	3648			
2	4753	1	3648			
2	4754	1	3648			
2	4755	1	3648			
2	4756	1	1606			
2	4757	1	1606			
2	4758	1	1606			
2	4759	1	1606			
2	4760	1	1606			
2	4761	1	3654			
2	4762	1	3654			
2	4763	1	3654			
2	4764	1	3654			
2	4765	1	1612			
2	4766	1	1612			
2	4767	1	1612			
2	4768	1	1615			
2	4769	1	1615			
2	4770	1	1615			
2	4771	1	1615			
2	4772	1	1619			
2	4773	1	1619			
2	4774	1	1619			
2	4775	1	1619			
2	4776	1	1619			
2	4777	1	1619			
2	4778	1	1619			
2	4779	1	1619			
2	4780	1	1624			
2	4781	1	1624			
2	4782	1	1624			
2	4783	1	1624			
2	4784	1	1624			
2	4785	1	1624			
2	4786	1	1624			
2	4787	1	1628			
2	4788	1	1628			
2	4789	1	1628			
2	4790	1	1628			
2	4791	1	1631			
2	4792	1	1631			
2	4793	1	1631			
2	4794	1	1631			
2	4795	1	1634			
2	4796	1	1634			
2	4797	1	1634			
2	4798	1	1634			
2	4799	1	1637			
2	4800	1	1637			
2	4801	1	1637			
2	4802	1	1637			
2	4803	1	1637			
2	4804	1	1642			
2	4805	1	1642			
2	4806	1	1642			
2	4807	1	1642			
2	4808	1	1642			
2	4809	1	1647			
2	4810	1	1647			
2	4811	1	1647			
2	4812	1	1647			
2	4813	1	1651			
2	4814	1	1651			
2	4815	1	1651			
2	4816	1	1651			
2	4817	1	1651			
2	4818	1	1656			
2	4819	1	1656			
2	4820	1	1656			
2	4821	1	1656			
2	4822	1	3723			
2	4823	1	3723			
2	4824	1	1676			
2	4825	1	1676			
2	4826	1	1676			
2	4827	1	1676			
2	4828	1	1676			
2	4829	1	1681			
2	4830	1	1681			
2	4831	1	1681			
2	4832	1	1681			
2	4833	1	1681			
2	4834	1	1686			
2	4835	1	1686			
2	4836	1	1686			
2	4837	1	1686			
2	4838	1	1686			
2	4839	1	1690			
2	4840	1	1690			
2	4841	1	1690			
2	4842	1	3737			
2	4843	1	3737			
2	4844	1	3754			
2	4845	1	3754			
2	4846	1	3754			
2	4847	1	1708			
2	4848	1	1708			
2	4849	1	3758			
2	4850	1	3758			
2	4851	1	3762			
2	4852	1	3762			
2	4853	1	3767			
2	4854	1	3767			
2	4855	1	3767			
2	4856	1	3771			
2	4857	1	3771			
2	4858	1	3775			
2	4859	1	3775			
2	4860	1	3608			
2	4861	1	3608			
2	4862	1	3608			
2	4863	1	1770			
2	4864	1	1770			
2	4865	1	1773			
2	4866	1	1773			
2	4867	1	3823			
2	4868	1	3823			
2	4869	1	3827			
2	4870	1	3827			
2	4871	1	3612			
2	4872	1	3612			
2	4873	1	3840			
2	4874	1	3840			
2	4875	1	1795			
2	4876	1	1795			
2	4877	1	3843			
2	4878	1	3843			
2	4879	1	1798			
2	4880	1	1798			
2	4881	1	3852			
2	4882	1	3852			
2	4883	1	3616			
2	4884	1	3616			
2	4885	1	3616			
2	4886	1	3616			
2	4887	1	3616			
2	4888	1	3864			
2	4889	1	3864			
2	4890	1	3870			
2	4891	1	3870			
2	4892	1	1827			
2	4893	1	1827			
2	4894	1	1833			
2	4895	1	1833			
2	4896	1	1833			
2	4897	1	1833			
2	4898	1	1836			
2	4899	1	1836			
2	4900	1	1836			
2	4901	1	1836			
2	4902	1	1836			
2	4903	1	1836			
2	4904	1	1841			
2	4905	1	1841			
2	4906	1	1841			
2	4907	1	1841			
2	4908	1	1841			
2	4909	1	1841			
2	4910	1	1841			
2	4911	1	1841			
2	4912	1	1841			
2	4913	1	1841			
2	4914	1	1885			
2	4915	1	1885			
2	4916	1	1888			
2	4917	1	1888			
2	4918	1	1894			
2	4919	1	1894			
2	4920	1	1897			
2	4921	1	1897			
2	4922	1	2046			
2	4923	1	2046			
