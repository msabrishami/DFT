1 0 0 6 0
1 1 0 4 0
1 2 0 3 0
1 3 0 8 0
1 4 0 2 0
1 5 0 6 0
1 6 0 5 0
1 7 0 8 0
1 8 0 3 0
1 9 0 3 0
1 10 0 8 0
1 11 0 3 0
1 12 0 1 0
1 13 0 1 0
1 14 0 1 0
1 15 0 4 0
1 16 0 4 0
1 17 0 1 0
1 18 0 1 0
1 19 0 1 0
1 20 0 1 0
1 21 0 1 0
1 22 0 1 0
1 23 0 4 0
1 24 0 4 0
1 25 0 4 0
1 26 0 4 0
1 27 0 4 0
1 28 0 4 0
1 29 0 4 0
1 30 0 3 0
1 31 0 4 0
1 32 0 2 0
1 33 0 4 0
1 34 0 2 0
1 35 0 2 0
1 36 0 2 0
1 37 0 1 0
1 38 0 2 0
1 39 0 2 0
1 40 0 5 0
1 41 0 5 0
1 42 0 5 0
1 43 0 5 0
1 44 0 5 0
1 45 0 5 0
1 46 0 5 0
1 47 0 5 0
1 48 0 2 0
1 49 0 8 0
1 50 0 8 0
1 51 0 8 0
1 52 0 8 0
1 53 0 8 0
1 54 0 3 0
1 55 0 1 0
1 56 0 1 0
1 57 0 5 0
1 58 0 1 0
1 59 0 1 0
3 60 5 0 1 96 
3 61 5 0 1 97 
3 62 5 0 1 98 
3 63 5 0 1 103 
3 64 5 0 1 139 
3 65 5 0 1 141 
3 66 5 0 1 148 
3 67 5 0 1 150 
3 68 5 0 1 151 
3 69 5 0 1 153 
3 70 5 0 1 164 
3 71 5 0 1 166 
3 72 5 0 1 168 
3 73 5 0 1 169 
3 74 5 0 1 170 
3 75 5 0 1 298 
3 76 5 0 1 299 
3 77 5 0 1 411 
3 78 5 0 1 425 
3 79 5 0 1 426 
3 80 5 0 1 427 
3 81 5 0 1 428 
3 82 5 0 1 436 
3 83 5 0 1 440 
3 84 5 0 1 441 
3 85 5 0 1 442 
0 86 6 1 4 443 449 453 456 
0 87 6 2 4 444 4 454 457 
0 88 7 2 3 464 470 475 
0 89 7 2 3 445 4 483 
0 90 6 1 4 446 450 484 458 
0 91 6 3 4 447 451 455 486 
0 92 6 1 4 489 476 497 12 
0 93 6 1 2 465 498 
0 94 6 1 3 490 499 14 
0 95 7 2 3 466 500 504 
0 96 7 1 3 467 501 477 
0 97 7 1 3 468 471 505 
0 98 7 1 3 469 472 478 
0 99 7 1 3 491 502 506 
0 100 7 1 3 492 503 479 
0 101 7 1 3 493 473 507 
0 102 7 1 3 494 474 480 
0 103 7 1 2 17 18 
0 104 3 2 2 19 20 
0 105 6 1 2 508 512 
0 106 3 1 2 509 513 
0 107 6 1 2 516 520 
0 108 3 1 2 517 521 
0 109 6 1 2 524 528 
0 110 3 1 2 525 529 
0 111 6 1 2 532 536 
0 112 3 1 2 533 537 
0 113 7 1 2 452 543 
0 114 5 5 1 59 
0 115 7 1 2 485 544 
0 116 7 1 2 459 545 
0 117 7 1 2 37 546 
0 118 6 2 2 495 39 
0 119 4 1 2 460 481 
0 120 7 1 2 461 482 
0 121 6 1 2 547 552 
0 122 3 1 2 548 553 
0 123 6 1 2 557 562 
0 124 3 1 2 558 563 
0 125 6 1 2 567 572 
0 126 3 1 2 568 573 
0 127 6 1 2 577 582 
0 128 3 1 2 578 583 
0 129 7 1 2 587 510 
0 130 7 1 2 588 514 
0 131 7 1 2 589 518 
0 132 7 1 2 590 522 
0 133 7 1 2 591 526 
0 134 7 1 2 627 55 
0 135 7 1 2 592 530 
0 136 7 1 2 628 56 
0 137 7 1 2 593 534 
0 138 7 1 2 629 58 
0 139 5 1 1 86 
0 140 5 1 1 637 
0 141 3 1 2 635 638 
0 142 5 1 1 639 
0 143 5 1 1 640 
0 144 5 1 1 90 
0 145 4 1 2 641 92 
0 146 3 1 2 642 93 
0 147 3 1 2 643 94 
0 148 5 1 1 99 
0 149 5 1 1 100 
0 150 5 1 1 101 
0 151 5 1 1 102 
0 152 6 1 2 21 646 
0 153 7 1 2 22 647 
0 154 6 2 2 105 106 
0 155 6 2 2 107 108 
0 156 6 2 2 109 110 
0 157 6 2 2 111 112 
0 158 5 5 1 648 
0 159 4 1 2 119 120 
0 160 6 2 2 121 122 
0 161 6 2 2 123 124 
0 162 6 2 2 125 126 
0 163 6 2 2 127 128 
0 164 3 1 2 636 140 
0 165 5 5 1 142 
0 166 5 1 1 143 
0 167 7 1 2 145 13 
0 168 5 1 1 146 
0 169 5 1 1 147 
0 170 5 1 1 152 
0 171 5 1 1 655 
0 172 5 1 1 657 
0 173 7 1 2 656 658 
0 174 5 1 1 659 
0 175 5 1 1 661 
0 176 7 1 2 660 662 
0 177 6 1 2 144 149 
0 178 5 1 1 668 
0 179 5 1 1 670 
0 180 7 1 2 669 671 
0 181 5 1 1 672 
0 182 5 1 1 674 
0 183 7 1 2 673 675 
0 184 7 1 2 594 663 
0 185 5 1 1 167 
0 186 7 1 2 171 172 
0 187 7 1 2 174 175 
0 188 7 4 3 653 676 487 
0 189 7 4 3 677 462 644 
0 190 6 4 3 678 645 488 
0 191 6 1 4 159 496 39 679 
0 192 6 1 3 680 654 463 
0 193 7 1 2 178 179 
0 194 7 1 2 181 182 
0 195 5 8 1 185 
0 196 4 2 2 173 186 
0 197 4 2 2 176 187 
0 198 6 8 2 191 177 
0 199 7 1 2 34 681 
0 200 7 1 2 649 685 
0 201 7 1 2 35 682 
0 202 7 1 2 650 686 
0 203 7 1 2 36 683 
0 204 7 1 2 651 687 
0 205 7 1 2 38 684 
0 206 7 1 2 652 688 
0 207 6 4 2 192 448 
0 208 3 1 2 664 689 
0 209 3 1 2 665 690 
0 210 3 1 2 666 691 
0 211 3 1 2 667 692 
0 212 4 2 2 180 193 
0 213 4 2 2 183 194 
0 214 6 1 2 539 701 
0 215 3 1 2 540 702 
0 216 6 1 2 703 32 
0 217 3 1 2 704 32 
0 218 7 1 2 511 705 
0 219 4 1 2 199 200 
0 220 7 1 2 515 706 
0 221 4 1 2 201 202 
0 222 7 1 2 519 707 
0 223 4 1 2 203 204 
0 224 7 1 2 523 708 
0 225 4 1 2 205 206 
0 226 7 1 2 34 713 
0 227 7 1 2 527 709 
0 228 7 1 2 35 714 
0 229 7 1 2 531 710 
0 230 7 1 2 36 715 
0 231 7 1 2 535 711 
0 232 7 1 2 38 716 
0 233 7 1 2 538 712 
0 234 6 1 2 541 717 
0 235 3 1 2 542 718 
0 236 6 1 2 719 48 
0 237 3 1 2 720 48 
0 238 7 1 2 693 549 
0 239 7 1 2 694 554 
0 240 7 1 2 695 559 
0 241 7 1 2 696 564 
0 242 7 1 2 697 569 
0 243 6 1 2 698 574 
0 244 6 1 2 699 579 
0 245 6 1 2 700 584 
0 246 6 2 2 214 215 
0 247 6 2 2 216 217 
0 248 4 1 2 113 218 
0 249 4 1 2 115 220 
0 250 4 1 2 116 222 
0 251 4 1 2 117 224 
0 252 4 1 2 226 227 
0 253 4 1 2 228 229 
0 254 4 1 2 230 231 
0 255 4 1 2 232 233 
0 256 6 2 2 234 235 
0 257 6 2 2 236 237 
0 258 5 1 1 721 
0 259 5 1 1 723 
0 260 7 1 2 722 724 
0 261 6 3 2 248 219 
0 262 6 3 2 249 221 
0 263 6 3 2 250 223 
0 264 6 3 2 251 225 
0 265 6 3 2 208 252 
0 266 6 3 2 209 253 
0 267 6 3 2 210 254 
0 268 6 3 2 211 255 
0 269 5 1 1 725 
0 270 5 1 1 727 
0 271 7 1 2 726 728 
0 272 7 1 2 258 259 
0 273 7 1 2 269 270 
0 274 6 2 2 729 550 
0 275 3 2 2 730 551 
0 276 7 1 2 619 731 
0 277 6 2 2 732 555 
0 278 3 4 2 733 556 
0 279 7 1 2 620 734 
0 280 6 2 2 735 560 
0 281 3 5 2 736 561 
0 282 7 1 2 621 737 
0 283 6 2 2 738 565 
0 284 3 4 2 739 566 
0 285 7 1 2 622 740 
0 286 6 2 2 741 570 
0 287 3 2 2 742 571 
0 288 7 1 2 623 743 
0 289 6 2 2 744 575 
0 290 3 4 2 745 576 
0 291 7 1 2 624 746 
0 292 6 2 2 747 580 
0 293 3 5 2 748 581 
0 294 7 1 2 625 749 
0 295 6 2 2 750 585 
0 296 3 4 2 751 586 
0 297 7 1 2 626 752 
0 298 4 1 2 260 272 
0 299 4 1 2 271 273 
0 300 5 2 1 753 
0 301 7 3 2 755 754 
0 302 4 1 2 276 238 
0 303 5 2 1 757 
0 304 7 3 2 759 758 
0 305 4 1 2 279 239 
0 306 5 3 1 763 
0 307 7 3 2 765 764 
0 308 4 1 2 282 240 
0 309 5 4 1 770 
0 310 7 3 2 772 771 
0 311 4 1 2 285 241 
0 312 5 2 1 776 
0 313 7 3 2 778 777 
0 314 4 1 2 288 242 
0 315 5 2 1 780 
0 316 7 3 2 782 781 
0 317 4 1 2 134 291 
0 318 5 3 1 786 
0 319 7 3 2 788 787 
0 320 4 1 2 136 294 
0 321 5 4 1 793 
0 322 7 3 2 795 794 
0 323 4 1 2 138 297 
0 324 6 1 2 796 630 
0 325 6 1 3 789 797 631 
0 326 6 1 4 783 790 798 632 
0 327 5 1 1 799 
0 328 7 1 2 603 801 
0 329 7 1 2 611 800 
0 330 5 1 1 804 
0 331 7 1 2 604 806 
0 332 7 1 2 612 805 
0 333 5 1 1 809 
0 334 7 1 2 605 812 
0 335 7 1 2 613 810 
0 336 5 1 1 815 
0 337 7 1 2 606 819 
0 338 7 1 2 614 816 
0 339 5 1 1 822 
0 340 7 1 2 607 824 
0 341 7 1 2 615 823 
0 342 5 1 1 827 
0 343 7 1 2 608 829 
0 344 7 1 2 616 828 
0 345 5 1 1 832 
0 346 7 1 2 609 835 
0 347 7 1 2 617 833 
0 348 5 1 1 838 
0 349 4 1 2 842 633 
0 350 7 1 2 843 634 
0 351 7 1 2 610 844 
0 352 7 1 2 618 839 
0 353 6 1 2 791 840 
0 354 6 1 2 784 834 
0 355 6 1 3 785 792 841 
0 356 6 1 2 766 817 
0 357 6 1 2 760 811 
0 358 6 1 3 761 767 818 
0 359 4 1 2 328 329 
0 360 4 1 2 331 332 
0 361 4 1 2 334 335 
0 362 4 1 2 337 338 
0 363 6 3 4 342 354 355 326 
0 364 4 1 2 340 341 
0 365 6 2 3 345 353 325 
0 366 4 1 2 343 344 
0 367 6 2 2 348 324 
0 368 4 1 2 346 347 
0 369 4 1 2 349 350 
0 370 4 1 2 351 352 
0 371 4 1 2 825 845 
0 372 7 1 2 826 846 
0 373 4 1 2 830 848 
0 374 7 1 2 831 849 
0 375 4 1 2 836 850 
0 376 7 1 2 837 851 
0 377 7 1 2 595 369 
0 378 6 1 2 779 847 
0 379 6 5 2 378 339 
0 380 4 1 2 371 372 
0 381 4 1 2 373 374 
0 382 4 1 2 375 376 
0 383 4 1 2 137 377 
0 384 4 1 2 820 852 
0 385 7 1 2 821 853 
0 386 7 1 2 596 380 
0 387 7 1 2 597 381 
0 388 7 1 2 598 382 
0 389 6 1 4 383 370 323 245 
0 390 6 1 2 773 854 
0 391 6 1 3 768 774 855 
0 392 6 1 4 762 769 775 856 
0 393 6 3 4 330 357 358 392 
0 394 6 2 3 333 356 391 
0 395 6 2 2 336 390 
0 396 4 1 2 384 385 
0 397 4 1 2 132 386 
0 398 4 1 2 133 387 
0 399 4 1 2 135 388 
0 400 5 1 1 389 
0 401 4 1 2 802 857 
0 402 7 1 2 803 858 
0 403 4 1 2 807 860 
0 404 7 1 2 808 861 
0 405 4 1 2 813 862 
0 406 7 1 2 814 863 
0 407 7 1 2 599 396 
0 408 6 1 3 397 364 314 
0 409 6 1 4 398 366 317 243 
0 410 6 1 4 399 368 320 244 
0 411 5 1 1 400 
0 412 6 1 2 859 756 
0 413 4 1 2 401 402 
0 414 4 1 2 403 404 
0 415 4 1 2 405 406 
0 416 4 1 2 131 407 
0 417 5 1 1 408 
0 418 5 1 1 409 
0 419 5 1 1 410 
0 420 7 1 2 327 412 
0 421 7 1 2 600 413 
0 422 7 1 2 601 414 
0 423 7 1 2 602 415 
0 424 6 1 3 416 362 311 
0 425 5 1 1 417 
0 426 5 1 1 418 
0 427 5 1 1 419 
0 428 5 1 1 420 
0 429 4 1 2 184 421 
0 430 4 1 2 129 422 
0 431 4 1 2 130 423 
0 432 5 1 1 424 
0 433 6 1 3 429 359 302 
0 434 6 1 3 430 360 305 
0 435 6 1 3 431 361 308 
0 436 5 1 1 432 
0 437 5 1 1 433 
0 438 5 1 1 434 
0 439 5 1 1 435 
0 440 5 1 1 437 
0 441 5 1 1 438 
0 442 5 1 1 439 
2 443 1 0
2 444 1 0
2 445 1 0
2 446 1 0
2 447 1 0
2 448 1 0
2 449 1 1
2 450 1 1
2 451 1 1
2 452 1 1
2 453 1 2
2 454 1 2
2 455 1 2
2 456 1 3
2 457 1 3
2 458 1 3
2 459 1 3
2 460 1 3
2 461 1 3
2 462 1 3
2 463 1 3
2 464 1 5
2 465 1 5
2 466 1 5
2 467 1 5
2 468 1 5
2 469 1 5
2 470 1 6
2 471 1 6
2 472 1 6
2 473 1 6
2 474 1 6
2 475 1 7
2 476 1 7
2 477 1 7
2 478 1 7
2 479 1 7
2 480 1 7
2 481 1 7
2 482 1 7
2 483 1 8
2 484 1 8
2 485 1 8
2 486 1 9
2 487 1 9
2 488 1 9
2 489 1 10
2 490 1 10
2 491 1 10
2 492 1 10
2 493 1 10
2 494 1 10
2 495 1 10
2 496 1 10
2 497 1 11
2 498 1 11
2 499 1 11
2 500 1 15
2 501 1 15
2 502 1 15
2 503 1 15
2 504 1 16
2 505 1 16
2 506 1 16
2 507 1 16
2 508 1 23
2 509 1 23
2 510 1 23
2 511 1 23
2 512 1 24
2 513 1 24
2 514 1 24
2 515 1 24
2 516 1 25
2 517 1 25
2 518 1 25
2 519 1 25
2 520 1 26
2 521 1 26
2 522 1 26
2 523 1 26
2 524 1 27
2 525 1 27
2 526 1 27
2 527 1 27
2 528 1 28
2 529 1 28
2 530 1 28
2 531 1 28
2 532 1 29
2 533 1 29
2 534 1 29
2 535 1 29
2 536 1 30
2 537 1 30
2 538 1 30
2 539 1 31
2 540 1 31
2 541 1 31
2 542 1 31
2 543 1 33
2 544 1 33
2 545 1 33
2 546 1 33
2 547 1 40
2 548 1 40
2 549 1 40
2 550 1 40
2 551 1 40
2 552 1 41
2 553 1 41
2 554 1 41
2 555 1 41
2 556 1 41
2 557 1 42
2 558 1 42
2 559 1 42
2 560 1 42
2 561 1 42
2 562 1 43
2 563 1 43
2 564 1 43
2 565 1 43
2 566 1 43
2 567 1 44
2 568 1 44
2 569 1 44
2 570 1 44
2 571 1 44
2 572 1 45
2 573 1 45
2 574 1 45
2 575 1 45
2 576 1 45
2 577 1 46
2 578 1 46
2 579 1 46
2 580 1 46
2 581 1 46
2 582 1 47
2 583 1 47
2 584 1 47
2 585 1 47
2 586 1 47
2 587 1 49
2 588 1 49
2 589 1 49
2 590 1 49
2 591 1 49
2 592 1 49
2 593 1 49
2 594 1 49
2 595 1 50
2 596 1 50
2 597 1 50
2 598 1 50
2 599 1 50
2 600 1 50
2 601 1 50
2 602 1 50
2 603 1 51
2 604 1 51
2 605 1 51
2 606 1 51
2 607 1 51
2 608 1 51
2 609 1 51
2 610 1 51
2 611 1 52
2 612 1 52
2 613 1 52
2 614 1 52
2 615 1 52
2 616 1 52
2 617 1 52
2 618 1 52
2 619 1 53
2 620 1 53
2 621 1 53
2 622 1 53
2 623 1 53
2 624 1 53
2 625 1 53
2 626 1 53
2 627 1 54
2 628 1 54
2 629 1 54
2 630 1 57
2 631 1 57
2 632 1 57
2 633 1 57
2 634 1 57
2 635 1 87
2 636 1 87
2 637 1 88
2 638 1 88
2 639 1 89
2 640 1 89
2 641 1 91
2 642 1 91
2 643 1 91
2 644 1 95
2 645 1 95
2 646 1 104
2 647 1 104
2 648 1 114
2 649 1 114
2 650 1 114
2 651 1 114
2 652 1 114
2 653 1 118
2 654 1 118
2 655 1 154
2 656 1 154
2 657 1 155
2 658 1 155
2 659 1 156
2 660 1 156
2 661 1 157
2 662 1 157
2 663 1 158
2 664 1 158
2 665 1 158
2 666 1 158
2 667 1 158
2 668 1 160
2 669 1 160
2 670 1 161
2 671 1 161
2 672 1 162
2 673 1 162
2 674 1 163
2 675 1 163
2 676 1 165
2 677 1 165
2 678 1 165
2 679 1 165
2 680 1 165
2 681 1 188
2 682 1 188
2 683 1 188
2 684 1 188
2 685 1 189
2 686 1 189
2 687 1 189
2 688 1 189
2 689 1 190
2 690 1 190
2 691 1 190
2 692 1 190
2 693 1 195
2 694 1 195
2 695 1 195
2 696 1 195
2 697 1 195
2 698 1 195
2 699 1 195
2 700 1 195
2 701 1 196
2 702 1 196
2 703 1 197
2 704 1 197
2 705 1 198
2 706 1 198
2 707 1 198
2 708 1 198
2 709 1 198
2 710 1 198
2 711 1 198
2 712 1 198
2 713 1 207
2 714 1 207
2 715 1 207
2 716 1 207
2 717 1 212
2 718 1 212
2 719 1 213
2 720 1 213
2 721 1 246
2 722 1 246
2 723 1 247
2 724 1 247
2 725 1 256
2 726 1 256
2 727 1 257
2 728 1 257
2 729 1 261
2 730 1 261
2 731 1 261
2 732 1 262
2 733 1 262
2 734 1 262
2 735 1 263
2 736 1 263
2 737 1 263
2 738 1 264
2 739 1 264
2 740 1 264
2 741 1 265
2 742 1 265
2 743 1 265
2 744 1 266
2 745 1 266
2 746 1 266
2 747 1 267
2 748 1 267
2 749 1 267
2 750 1 268
2 751 1 268
2 752 1 268
2 753 1 274
2 754 1 274
2 755 1 275
2 756 1 275
2 757 1 277
2 758 1 277
2 759 1 278
2 760 1 278
2 761 1 278
2 762 1 278
2 763 1 280
2 764 1 280
2 765 1 281
2 766 1 281
2 767 1 281
2 768 1 281
2 769 1 281
2 770 1 283
2 771 1 283
2 772 1 284
2 773 1 284
2 774 1 284
2 775 1 284
2 776 1 286
2 777 1 286
2 778 1 287
2 779 1 287
2 780 1 289
2 781 1 289
2 782 1 290
2 783 1 290
2 784 1 290
2 785 1 290
2 786 1 292
2 787 1 292
2 788 1 293
2 789 1 293
2 790 1 293
2 791 1 293
2 792 1 293
2 793 1 295
2 794 1 295
2 795 1 296
2 796 1 296
2 797 1 296
2 798 1 296
2 799 1 300
2 800 1 300
2 801 1 301
2 802 1 301
2 803 1 301
2 804 1 303
2 805 1 303
2 806 1 304
2 807 1 304
2 808 1 304
2 809 1 306
2 810 1 306
2 811 1 306
2 812 1 307
2 813 1 307
2 814 1 307
2 815 1 309
2 816 1 309
2 817 1 309
2 818 1 309
2 819 1 310
2 820 1 310
2 821 1 310
2 822 1 312
2 823 1 312
2 824 1 313
2 825 1 313
2 826 1 313
2 827 1 315
2 828 1 315
2 829 1 316
2 830 1 316
2 831 1 316
2 832 1 318
2 833 1 318
2 834 1 318
2 835 1 319
2 836 1 319
2 837 1 319
2 838 1 321
2 839 1 321
2 840 1 321
2 841 1 321
2 842 1 322
2 843 1 322
2 844 1 322
2 845 1 363
2 846 1 363
2 847 1 363
2 848 1 365
2 849 1 365
2 850 1 367
2 851 1 367
2 852 1 379
2 853 1 379
2 854 1 379
2 855 1 379
2 856 1 379
2 857 1 393
2 858 1 393
2 859 1 393
2 860 1 394
2 861 1 394
2 862 1 395
2 863 1 395
