1 N1 0 7 0
1 N8 0 7 0
1 N15 0 7 0
1 N22 0 7 0
1 N29 0 7 0
1 N36 0 7 0
1 N43 0 7 0
1 N50 0 7 0
1 N57 0 7 0
1 N64 0 7 0
1 N71 0 7 0
1 N78 0 7 0
1 N85 0 7 0
1 N92 0 7 0
1 N99 0 7 0
1 N106 0 7 0
1 N113 0 7 0
1 N120 0 7 0
1 N127 0 7 0
1 N134 0 7 0
1 N141 0 7 0
1 N148 0 7 0
1 N155 0 7 0
1 N162 0 7 0
1 N169 0 7 0
1 N176 0 7 0
1 N183 0 7 0
1 N190 0 7 0
1 N197 0 7 0
1 N204 0 7 0
1 N211 0 7 0
1 N218 0 7 0
1 N225 0 3 0
1 N226 0 3 0
1 N227 0 3 0
1 N228 0 3 0
1 N229 0 3 0
1 N230 0 3 0
1 N231 0 3 0
1 N232 0 2 0
1 N233 0 17 0
2 N1-1 1 N1 
2 N1-2 1 N1 
2 N1-3 1 N1 
2 N1-4 1 N1 
2 N1-5 1 N1 
2 N1-6 1 N1 
2 N1-7 1 N1 
2 N8-1 1 N8 
2 N8-2 1 N8 
2 N8-3 1 N8 
2 N8-4 1 N8 
2 N8-5 1 N8 
2 N8-6 1 N8 
2 N8-7 1 N8 
2 N15-1 1 N15 
2 N15-2 1 N15 
2 N15-3 1 N15 
2 N15-4 1 N15 
2 N15-5 1 N15 
2 N15-6 1 N15 
2 N15-7 1 N15 
2 N22-1 1 N22 
2 N22-2 1 N22 
2 N22-3 1 N22 
2 N22-4 1 N22 
2 N22-5 1 N22 
2 N22-6 1 N22 
2 N22-7 1 N22 
2 N29-1 1 N29 
2 N29-2 1 N29 
2 N29-3 1 N29 
2 N29-4 1 N29 
2 N29-5 1 N29 
2 N29-6 1 N29 
2 N29-7 1 N29 
2 N36-1 1 N36 
2 N36-2 1 N36 
2 N36-3 1 N36 
2 N36-4 1 N36 
2 N36-5 1 N36 
2 N36-6 1 N36 
2 N36-7 1 N36 
2 N43-1 1 N43 
2 N43-2 1 N43 
2 N43-3 1 N43 
2 N43-4 1 N43 
2 N43-5 1 N43 
2 N43-6 1 N43 
2 N43-7 1 N43 
2 N50-1 1 N50 
2 N50-2 1 N50 
2 N50-3 1 N50 
2 N50-4 1 N50 
2 N50-5 1 N50 
2 N50-6 1 N50 
2 N50-7 1 N50 
2 N57-1 1 N57 
2 N57-2 1 N57 
2 N57-3 1 N57 
2 N57-4 1 N57 
2 N57-5 1 N57 
2 N57-6 1 N57 
2 N57-7 1 N57 
2 N64-1 1 N64 
2 N64-2 1 N64 
2 N64-3 1 N64 
2 N64-4 1 N64 
2 N64-5 1 N64 
2 N64-6 1 N64 
2 N64-7 1 N64 
2 N71-1 1 N71 
2 N71-2 1 N71 
2 N71-3 1 N71 
2 N71-4 1 N71 
2 N71-5 1 N71 
2 N71-6 1 N71 
2 N71-7 1 N71 
2 N78-1 1 N78 
2 N78-2 1 N78 
2 N78-3 1 N78 
2 N78-4 1 N78 
2 N78-5 1 N78 
2 N78-6 1 N78 
2 N78-7 1 N78 
2 N85-1 1 N85 
2 N85-2 1 N85 
2 N85-3 1 N85 
2 N85-4 1 N85 
2 N85-5 1 N85 
2 N85-6 1 N85 
2 N85-7 1 N85 
2 N92-1 1 N92 
2 N92-2 1 N92 
2 N92-3 1 N92 
2 N92-4 1 N92 
2 N92-5 1 N92 
2 N92-6 1 N92 
2 N92-7 1 N92 
2 N99-1 1 N99 
2 N99-2 1 N99 
2 N99-3 1 N99 
2 N99-4 1 N99 
2 N99-5 1 N99 
2 N99-6 1 N99 
2 N99-7 1 N99 
2 N106-1 1 N106 
2 N106-2 1 N106 
2 N106-3 1 N106 
2 N106-4 1 N106 
2 N106-5 1 N106 
2 N106-6 1 N106 
2 N106-7 1 N106 
2 N113-1 1 N113 
2 N113-2 1 N113 
2 N113-3 1 N113 
2 N113-4 1 N113 
2 N113-5 1 N113 
2 N113-6 1 N113 
2 N113-7 1 N113 
2 N120-1 1 N120 
2 N120-2 1 N120 
2 N120-3 1 N120 
2 N120-4 1 N120 
2 N120-5 1 N120 
2 N120-6 1 N120 
2 N120-7 1 N120 
2 N127-1 1 N127 
2 N127-2 1 N127 
2 N127-3 1 N127 
2 N127-4 1 N127 
2 N127-5 1 N127 
2 N127-6 1 N127 
2 N127-7 1 N127 
2 N134-1 1 N134 
2 N134-2 1 N134 
2 N134-3 1 N134 
2 N134-4 1 N134 
2 N134-5 1 N134 
2 N134-6 1 N134 
2 N134-7 1 N134 
2 N141-1 1 N141 
2 N141-2 1 N141 
2 N141-3 1 N141 
2 N141-4 1 N141 
2 N141-5 1 N141 
2 N141-6 1 N141 
2 N141-7 1 N141 
2 N148-1 1 N148 
2 N148-2 1 N148 
2 N148-3 1 N148 
2 N148-4 1 N148 
2 N148-5 1 N148 
2 N148-6 1 N148 
2 N148-7 1 N148 
2 N155-1 1 N155 
2 N155-2 1 N155 
2 N155-3 1 N155 
2 N155-4 1 N155 
2 N155-5 1 N155 
2 N155-6 1 N155 
2 N155-7 1 N155 
2 N162-1 1 N162 
2 N162-2 1 N162 
2 N162-3 1 N162 
2 N162-4 1 N162 
2 N162-5 1 N162 
2 N162-6 1 N162 
2 N162-7 1 N162 
2 N169-1 1 N169 
2 N169-2 1 N169 
2 N169-3 1 N169 
2 N169-4 1 N169 
2 N169-5 1 N169 
2 N169-6 1 N169 
2 N169-7 1 N169 
2 N176-1 1 N176 
2 N176-2 1 N176 
2 N176-3 1 N176 
2 N176-4 1 N176 
2 N176-5 1 N176 
2 N176-6 1 N176 
2 N176-7 1 N176 
2 N183-1 1 N183 
2 N183-2 1 N183 
2 N183-3 1 N183 
2 N183-4 1 N183 
2 N183-5 1 N183 
2 N183-6 1 N183 
2 N183-7 1 N183 
2 N190-1 1 N190 
2 N190-2 1 N190 
2 N190-3 1 N190 
2 N190-4 1 N190 
2 N190-5 1 N190 
2 N190-6 1 N190 
2 N190-7 1 N190 
2 N197-1 1 N197 
2 N197-2 1 N197 
2 N197-3 1 N197 
2 N197-4 1 N197 
2 N197-5 1 N197 
2 N197-6 1 N197 
2 N197-7 1 N197 
2 N204-1 1 N204 
2 N204-2 1 N204 
2 N204-3 1 N204 
2 N204-4 1 N204 
2 N204-5 1 N204 
2 N204-6 1 N204 
2 N204-7 1 N204 
2 N211-1 1 N211 
2 N211-2 1 N211 
2 N211-3 1 N211 
2 N211-4 1 N211 
2 N211-5 1 N211 
2 N211-6 1 N211 
2 N211-7 1 N211 
2 N218-1 1 N218 
2 N218-2 1 N218 
2 N218-3 1 N218 
2 N218-4 1 N218 
2 N218-5 1 N218 
2 N218-6 1 N218 
2 N218-7 1 N218 
2 N225-1 1 N225 
2 N225-2 1 N225 
2 N225-3 1 N225 
2 N226-1 1 N226 
2 N226-2 1 N226 
2 N226-3 1 N226 
2 N227-1 1 N227 
2 N227-2 1 N227 
2 N227-3 1 N227 
2 N228-1 1 N228 
2 N228-2 1 N228 
2 N228-3 1 N228 
2 N229-1 1 N229 
2 N229-2 1 N229 
2 N229-3 1 N229 
2 N230-1 1 N230 
2 N230-2 1 N230 
2 N230-3 1 N230 
2 N231-1 1 N231 
2 N231-2 1 N231 
2 N231-3 1 N231 
2 N232-1 1 N232 
2 N232-2 1 N232 
2 N233-1 1 N233 
2 N233-2 1 N233 
2 N233-3 1 N233 
2 N233-4 1 N233 
2 N233-5 1 N233 
2 N233-6 1 N233 
2 N233-7 1 N233 
2 N233-8 1 N233 
2 N233-9 1 N233 
2 N233-10 1 N233 
2 N233-11 1 N233 
2 N233-12 1 N233 
2 N233-13 1 N233 
2 N233-14 1 N233 
2 N233-15 1 N233 
2 N233-16 1 N233 
2 N233-17 1 N233 
0 n640 5 2 1 N232-1
0 n648 6 1 2 N232-2 N233-2
0 n679 7 1 2 N230-1 N233-3
0 n687 6 1 2 N230-3 N233-4
0 n739 7 1 2 N228-1 N233-5
0 n747 6 1 2 N228-3 N233-6
0 n702 5 4 1 N106-6
0 n777 7 1 2 N227-1 N233-7
0 n785 6 1 2 N227-3 N233-8
0 n699 5 4 1 N99-7
0 n815 7 1 2 N226-1 N233-9
0 n823 6 1 2 N226-3 N233-10
0 n715 5 4 1 N204-7
0 n660 5 4 1 N218-7
0 n659 5 4 1 N190-7
0 n714 5 4 1 N176-7
0 n698 5 4 1 N92-7
0 n881 7 1 2 N225-1 N233-11
0 n889 6 1 2 N225-3 N233-12
0 n718 5 4 1 N120-7
0 n663 5 4 1 N134-7
0 n719 5 4 1 N148-7
0 n664 5 4 1 N162-7
0 n703 5 4 1 N85-7
0 n947 7 1 2 N229-1 N233-13
0 n955 6 1 2 N229-3 N233-14
0 n932 5 4 1 N29-6
0 n865 5 4 1 N36-7
0 n800 5 4 1 N43-6
0 n758 5 4 1 N50-7
0 n901 5 4 1 N113-6
0 n917 5 4 1 N141-7
0 n848 5 4 1 N169-6
0 n835 5 4 1 N197-7
0 n994 7 1 2 N231-1 N233-15
0 n641 5 8 1 N233-16
0 n1002 6 1 2 N231-3 N233-17
0 n931 5 4 1 N1-6
0 n799 5 4 1 N15-7
0 n762 5 4 1 N22-6
0 n862 5 4 1 N8-7
0 n796 5 4 1 N71-6
0 n759 5 4 1 N78-7
0 n928 5 4 1 N57-6
0 n866 5 4 1 N64-7
0 n898 5 4 1 N127-6
0 n914 5 4 1 N155-7
0 n851 5 4 1 N183-6
0 n832 5 4 1 N211-7
2 n640-1 1 n640 
2 n640-2 1 n640 
2 n702-1 1 n702 
2 n702-2 1 n702 
2 n702-3 1 n702 
2 n702-4 1 n702 
2 n699-1 1 n699 
2 n699-2 1 n699 
2 n699-3 1 n699 
2 n699-4 1 n699 
2 n715-1 1 n715 
2 n715-2 1 n715 
2 n715-3 1 n715 
2 n715-4 1 n715 
2 n660-1 1 n660 
2 n660-2 1 n660 
2 n660-3 1 n660 
2 n660-4 1 n660 
2 n659-1 1 n659 
2 n659-2 1 n659 
2 n659-3 1 n659 
2 n659-4 1 n659 
2 n714-1 1 n714 
2 n714-2 1 n714 
2 n714-3 1 n714 
2 n714-4 1 n714 
2 n698-1 1 n698 
2 n698-2 1 n698 
2 n698-3 1 n698 
2 n698-4 1 n698 
2 n718-1 1 n718 
2 n718-2 1 n718 
2 n718-3 1 n718 
2 n718-4 1 n718 
2 n663-1 1 n663 
2 n663-2 1 n663 
2 n663-3 1 n663 
2 n663-4 1 n663 
2 n719-1 1 n719 
2 n719-2 1 n719 
2 n719-3 1 n719 
2 n719-4 1 n719 
2 n664-1 1 n664 
2 n664-2 1 n664 
2 n664-3 1 n664 
2 n664-4 1 n664 
2 n703-1 1 n703 
2 n703-2 1 n703 
2 n703-3 1 n703 
2 n703-4 1 n703 
2 n932-1 1 n932 
2 n932-2 1 n932 
2 n932-3 1 n932 
2 n932-4 1 n932 
2 n865-1 1 n865 
2 n865-2 1 n865 
2 n865-3 1 n865 
2 n865-4 1 n865 
2 n800-1 1 n800 
2 n800-2 1 n800 
2 n800-3 1 n800 
2 n800-4 1 n800 
2 n758-1 1 n758 
2 n758-2 1 n758 
2 n758-3 1 n758 
2 n758-4 1 n758 
2 n901-1 1 n901 
2 n901-2 1 n901 
2 n901-3 1 n901 
2 n901-4 1 n901 
2 n917-1 1 n917 
2 n917-2 1 n917 
2 n917-3 1 n917 
2 n917-4 1 n917 
2 n848-1 1 n848 
2 n848-2 1 n848 
2 n848-3 1 n848 
2 n848-4 1 n848 
2 n835-1 1 n835 
2 n835-2 1 n835 
2 n835-3 1 n835 
2 n835-4 1 n835 
2 n641-1 1 n641 
2 n641-2 1 n641 
2 n641-3 1 n641 
2 n641-4 1 n641 
2 n641-5 1 n641 
2 n641-6 1 n641 
2 n641-7 1 n641 
2 n641-8 1 n641 
2 n931-1 1 n931 
2 n931-2 1 n931 
2 n931-3 1 n931 
2 n931-4 1 n931 
2 n799-1 1 n799 
2 n799-2 1 n799 
2 n799-3 1 n799 
2 n799-4 1 n799 
2 n762-1 1 n762 
2 n762-2 1 n762 
2 n762-3 1 n762 
2 n762-4 1 n762 
2 n862-1 1 n862 
2 n862-2 1 n862 
2 n862-3 1 n862 
2 n862-4 1 n862 
2 n796-1 1 n796 
2 n796-2 1 n796 
2 n796-3 1 n796 
2 n796-4 1 n796 
2 n759-1 1 n759 
2 n759-2 1 n759 
2 n759-3 1 n759 
2 n759-4 1 n759 
2 n928-1 1 n928 
2 n928-2 1 n928 
2 n928-3 1 n928 
2 n928-4 1 n928 
2 n866-1 1 n866 
2 n866-2 1 n866 
2 n866-3 1 n866 
2 n866-4 1 n866 
2 n898-1 1 n898 
2 n898-2 1 n898 
2 n898-3 1 n898 
2 n898-4 1 n898 
2 n914-1 1 n914 
2 n914-2 1 n914 
2 n914-3 1 n914 
2 n914-4 1 n914 
2 n851-1 1 n851 
2 n851-2 1 n851 
2 n851-3 1 n851 
2 n851-4 1 n851 
2 n832-1 1 n832 
2 n832-2 1 n832 
2 n832-3 1 n832 
2 n832-4 1 n832 
0 n638 4 1 2 n640-1 n641-1
0 n658 6 1 2 N218-3 n659-1
0 n657 6 1 2 N190-3 n660-1
0 n662 4 1 2 N162-3 n663-1
0 n661 4 1 2 N134-3 n664-1
0 n668 6 1 2 N162-4 n663-2
0 n667 6 1 2 N134-4 n664-2
0 n670 4 1 2 N218-4 n659-2
0 n669 4 1 2 N190-4 n660-2
0 n697 6 1 2 N99-3 n698-1
0 n696 6 1 2 N92-3 n699-1
0 n701 4 1 2 N85-3 n702-1
0 n700 4 1 2 N106-3 n703-1
0 n707 6 1 2 N85-4 n702-2
0 n706 6 1 2 N106-4 n703-2
0 n709 4 1 2 N99-4 n698-2
0 n708 4 1 2 N92-4 n699-2
0 n713 6 1 2 N204-3 n714-1
0 n712 6 1 2 N176-3 n715-1
0 n717 4 1 2 N148-3 n718-1
0 n716 4 1 2 N120-3 n719-1
0 n723 6 1 2 N148-4 n718-2
0 n722 6 1 2 N120-4 n719-2
0 n725 4 1 2 N204-4 n714-2
0 n724 4 1 2 N176-4 n715-2
0 n757 6 1 2 N78-3 n758-1
0 n756 6 1 2 N50-3 n759-1
0 n761 4 1 2 N22-3 n702-3
0 n760 4 1 2 N106-5 n762-1
0 n766 6 1 2 N22-4 n702-4
0 n765 6 1 2 N106-7 n762-2
0 n768 4 1 2 N78-4 n758-2
0 n767 4 1 2 N50-4 n759-2
0 n795 6 1 2 N99-5 n796-1
0 n794 6 1 2 N71-3 n699-3
0 n798 4 1 2 N43-3 n799-1
0 n797 4 1 2 N15-3 n800-1
0 n804 6 1 2 N43-4 n799-2
0 n803 6 1 2 N15-4 n800-2
0 n806 4 1 2 N99-6 n796-2
0 n805 4 1 2 N71-4 n699-4
0 n831 6 1 2 N218-5 n832-1
0 n830 6 1 2 N211-3 n660-3
0 n834 4 1 2 N204-5 n835-1
0 n833 4 1 2 N197-3 n715-3
0 n839 6 1 2 N204-6 n835-2
0 n838 6 1 2 N197-4 n715-4
0 n841 4 1 2 N218-6 n832-2
0 n840 4 1 2 N211-4 n660-4
0 n847 6 1 2 N176-5 n848-1
0 n846 6 1 2 N169-3 n714-3
0 n850 4 1 2 N190-5 n851-1
0 n849 4 1 2 N183-3 n659-3
0 n855 6 1 2 N190-6 n851-2
0 n854 6 1 2 N183-4 n659-4
0 n857 4 1 2 N176-6 n848-2
0 n856 4 1 2 N169-4 n714-4
0 n861 6 1 2 N92-5 n862-1
0 n860 6 1 2 N8-3 n698-3
0 n864 4 1 2 N64-3 n865-1
0 n863 4 1 2 N36-3 n866-1
0 n870 6 1 2 N64-4 n865-2
0 n869 6 1 2 N36-4 n866-2
0 n872 4 1 2 N92-6 n862-2
0 n871 4 1 2 N8-4 n698-4
0 n897 6 1 2 N134-5 n898-1
0 n896 6 1 2 N127-3 n663-3
0 n900 4 1 2 N120-5 n901-1
0 n899 4 1 2 N113-3 n718-3
0 n905 6 1 2 N120-6 n901-2
0 n904 6 1 2 N113-4 n718-4
0 n907 4 1 2 N134-6 n898-2
0 n906 4 1 2 N127-4 n663-4
0 n913 6 1 2 N162-5 n914-1
0 n912 6 1 2 N155-3 n664-3
0 n916 4 1 2 N148-5 n917-1
0 n915 4 1 2 N141-3 n719-3
0 n921 6 1 2 N148-6 n917-2
0 n920 6 1 2 N141-4 n719-4
0 n923 4 1 2 N162-6 n914-2
0 n922 4 1 2 N155-4 n664-4
0 n927 6 1 2 N85-5 n928-1
0 n926 6 1 2 N57-3 n703-3
0 n930 4 1 2 N29-3 n931-1
0 n929 4 1 2 N1-3 n932-1
0 n936 6 1 2 N29-4 n931-2
0 n935 6 1 2 N1-4 n932-2
0 n938 4 1 2 N85-6 n928-2
0 n937 4 1 2 N57-4 n703-4
0 n965 6 1 2 N50-5 n800-3
0 n964 6 1 2 N43-5 n758-3
0 n967 4 1 2 N36-5 n932-3
0 n966 4 1 2 N29-5 n865-3
0 n971 6 1 2 N36-6 n932-4
0 n970 6 1 2 N29-7 n865-4
0 n973 4 1 2 N50-6 n800-4
0 n972 4 1 2 N43-7 n758-4
0 n977 6 1 2 N197-5 n848-3
0 n976 6 1 2 N169-5 n835-3
0 n979 4 1 2 N141-5 n901-3
0 n978 4 1 2 N113-5 n917-3
0 n983 6 1 2 N141-6 n901-4
0 n982 6 1 2 N113-7 n917-4
0 n985 4 1 2 N197-6 n848-4
0 n984 4 1 2 N169-7 n835-4
0 n1010 6 1 2 N8-5 n762-3
0 n1009 6 1 2 N22-5 n862-3
0 n1012 4 1 2 N15-5 n931-3
0 n1011 4 1 2 N1-5 n799-3
0 n1016 6 1 2 N15-6 n931-4
0 n1015 6 1 2 N1-7 n799-4
0 n1018 4 1 2 N8-6 n762-4
0 n1017 4 1 2 N22-7 n862-4
0 n1024 6 1 2 N64-5 n928-3
0 n1023 6 1 2 N57-5 n866-3
0 n1026 4 1 2 N78-5 n796-3
0 n1025 4 1 2 N71-5 n759-3
0 n1030 6 1 2 N78-6 n796-4
0 n1029 6 1 2 N71-7 n759-4
0 n1032 4 1 2 N64-6 n928-4
0 n1031 4 1 2 N57-7 n866-4
0 n1036 6 1 2 N211-5 n851-3
0 n1035 6 1 2 N183-5 n832-3
0 n1038 4 1 2 N155-5 n898-3
0 n1037 4 1 2 N127-5 n914-3
0 n1042 6 1 2 N155-6 n898-4
0 n1041 6 1 2 N127-7 n914-4
0 n1044 4 1 2 N211-6 n851-4
0 n1043 4 1 2 N183-7 n832-4
0 n656 6 1 2 n657 n658
0 n655 4 1 2 n661 n662
0 n666 6 1 2 n667 n668
0 n665 4 1 2 n669 n670
0 n695 6 1 2 n696 n697
0 n694 4 1 2 n700 n701
0 n705 6 1 2 n706 n707
0 n704 4 1 2 n708 n709
0 n711 6 1 2 n712 n713
0 n710 4 1 2 n716 n717
0 n721 6 1 2 n722 n723
0 n720 4 1 2 n724 n725
0 n755 6 1 2 n756 n757
0 n754 4 1 2 n760 n761
0 n764 6 1 2 n765 n766
0 n763 4 1 2 n767 n768
0 n793 6 1 2 n794 n795
0 n792 4 1 2 n797 n798
0 n802 6 1 2 n803 n804
0 n801 4 1 2 n805 n806
0 n829 6 1 2 n830 n831
0 n828 4 1 2 n833 n834
0 n837 6 1 2 n838 n839
0 n836 4 1 2 n840 n841
0 n845 6 1 2 n846 n847
0 n844 4 1 2 n849 n850
0 n853 6 1 2 n854 n855
0 n852 4 1 2 n856 n857
0 n859 6 1 2 n860 n861
0 n858 4 1 2 n863 n864
0 n868 6 1 2 n869 n870
0 n867 4 1 2 n871 n872
0 n895 6 1 2 n896 n897
0 n894 4 1 2 n899 n900
0 n903 6 1 2 n904 n905
0 n902 4 1 2 n906 n907
0 n911 6 1 2 n912 n913
0 n910 4 1 2 n915 n916
0 n919 6 1 2 n920 n921
0 n918 4 1 2 n922 n923
0 n925 6 1 2 n926 n927
0 n924 4 1 2 n929 n930
0 n934 6 1 2 n935 n936
0 n933 4 1 2 n937 n938
0 n963 6 1 2 n964 n965
0 n962 4 1 2 n966 n967
0 n969 6 1 2 n970 n971
0 n968 4 1 2 n972 n973
0 n975 6 1 2 n976 n977
0 n974 4 1 2 n978 n979
0 n981 6 1 2 n982 n983
0 n980 4 1 2 n984 n985
0 n1008 6 1 2 n1009 n1010
0 n1007 4 1 2 n1011 n1012
0 n1014 6 1 2 n1015 n1016
0 n1013 4 1 2 n1017 n1018
0 n1022 6 1 2 n1023 n1024
0 n1021 4 1 2 n1025 n1026
0 n1028 6 1 2 n1029 n1030
0 n1027 4 1 2 n1031 n1032
0 n1034 6 1 2 n1035 n1036
0 n1033 4 1 2 n1037 n1038
0 n1040 6 1 2 n1041 n1042
0 n1039 4 1 2 n1043 n1044
0 n634 6 2 2 n655 n656
0 n635 6 2 2 n665 n666
0 n693 6 1 2 n694 n695
0 n692 6 1 2 n704 n705
0 n675 6 2 2 n710 n711
0 n676 6 2 2 n720 n721
0 n735 6 2 2 n754 n755
0 n736 6 2 2 n763 n764
0 n773 6 2 2 n792 n793
0 n774 6 2 2 n801 n802
0 n827 6 1 2 n828 n829
0 n826 6 1 2 n836 n837
0 n843 6 1 2 n844 n845
0 n842 6 1 2 n852 n853
0 n811 6 2 2 n858 n859
0 n812 6 2 2 n867 n868
0 n893 6 1 2 n894 n895
0 n892 6 1 2 n902 n903
0 n909 6 1 2 n910 n911
0 n908 6 1 2 n918 n919
0 n877 6 2 2 n924 n925
0 n878 6 2 2 n933 n934
0 n961 6 1 2 n962 n963
0 n960 6 1 2 n968 n969
0 n943 6 2 2 n974 n975
0 n944 6 2 2 n980 n981
0 n1006 6 1 2 n1007 n1008
0 n1005 6 1 2 n1013 n1014
0 n1020 6 1 2 n1021 n1022
0 n1019 6 1 2 n1027 n1028
0 n990 6 2 2 n1033 n1034
0 n991 6 2 2 n1039 n1040
0 n652 6 3 2 n692 n693
0 n751 6 3 2 n826 n827
0 n789 6 3 2 n842 n843
0 n791 6 3 2 n892 n893
0 n753 6 3 2 n908 n909
0 n654 6 3 2 n960 n961
0 n958 6 3 2 n1005 n1006
0 n690 6 3 2 n1019 n1020
2 n634-1 1 n634 
2 n634-2 1 n634 
2 n635-1 1 n635 
2 n635-2 1 n635 
2 n675-1 1 n675 
2 n675-2 1 n675 
2 n676-1 1 n676 
2 n676-2 1 n676 
2 n735-1 1 n735 
2 n735-2 1 n735 
2 n736-1 1 n736 
2 n736-2 1 n736 
2 n773-1 1 n773 
2 n773-2 1 n773 
2 n774-1 1 n774 
2 n774-2 1 n774 
2 n811-1 1 n811 
2 n811-2 1 n811 
2 n812-1 1 n812 
2 n812-2 1 n812 
2 n877-1 1 n877 
2 n877-2 1 n877 
2 n878-1 1 n878 
2 n878-2 1 n878 
2 n943-1 1 n943 
2 n943-2 1 n943 
2 n944-1 1 n944 
2 n944-2 1 n944 
2 n990-1 1 n990 
2 n990-2 1 n990 
2 n991-1 1 n991 
2 n991-2 1 n991 
0 n633 6 1 2 n634-1 n635-1
0 n643 7 1 2 n634-2 n635-2
0 n674 6 1 2 n675-1 n676-1
0 n682 7 1 2 n675-2 n676-2
0 n734 6 1 2 n735-1 n736-1
0 n742 7 1 2 n735-2 n736-2
0 n772 6 1 2 n773-1 n774-1
0 n780 7 1 2 n773-2 n774-2
0 n810 6 1 2 n811-1 n812-1
0 n818 7 1 2 n811-2 n812-2
0 n876 6 1 2 n877-1 n878-1
0 n884 7 1 2 n877-2 n878-2
0 n942 6 1 2 n943-1 n944-1
0 n950 7 1 2 n943-2 n944-2
0 n989 6 1 2 n990-1 n991-1
0 n997 7 1 2 n990-2 n991-2
2 n652-1 1 n652 
2 n652-2 1 n652 
2 n652-3 1 n652 
2 n751-1 1 n751 
2 n751-2 1 n751 
2 n751-3 1 n751 
2 n789-1 1 n789 
2 n789-2 1 n789 
2 n789-3 1 n789 
2 n791-1 1 n791 
2 n791-2 1 n791 
2 n791-3 1 n791 
2 n753-1 1 n753 
2 n753-2 1 n753 
2 n753-3 1 n753 
2 n654-1 1 n654 
2 n654-2 1 n654 
2 n654-3 1 n654 
2 n958-1 1 n958 
2 n958-2 1 n958 
2 n958-3 1 n958 
2 n690-1 1 n690 
2 n690-2 1 n690 
2 n690-3 1 n690 
0 n653 5 2 1 n652-2
0 n752 5 2 1 n751-2
0 n790 5 2 1 n789-3
0 n788 5 2 1 n791-2
0 n750 5 2 1 n753-3
0 n651 5 2 1 n654-2
0 n959 5 2 1 n958-2
0 n691 5 2 1 n690-3
2 n653-1 1 n653 
2 n653-2 1 n653 
2 n752-1 1 n752 
2 n752-2 1 n752 
2 n790-1 1 n790 
2 n790-2 1 n790 
2 n788-1 1 n788 
2 n788-2 1 n788 
2 n750-1 1 n750 
2 n750-2 1 n750 
2 n651-1 1 n651 
2 n651-2 1 n651 
2 n959-1 1 n959 
2 n959-2 1 n959 
2 n691-1 1 n691 
2 n691-2 1 n691 
0 n650 6 1 2 n652-1 n651-1
0 n649 6 1 2 n653-1 n654-1
0 n689 6 1 2 n653-2 n690-1
0 n688 6 1 2 n652-3 n691-1
0 n749 6 1 2 n751-1 n750-1
0 n748 6 1 2 n752-1 n753-1
0 n787 6 1 2 n789-1 n788-1
0 n786 6 1 2 n790-1 n791-1
0 n825 6 1 2 n752-2 n789-2
0 n824 6 1 2 n751-3 n790-2
0 n891 6 1 2 n788-2 n753-2
0 n890 6 1 2 n791-3 n750-2
0 n957 6 1 2 n651-2 n958-1
0 n956 6 1 2 n654-3 n959-1
0 n1004 6 1 2 n959-2 n690-2
0 n1003 6 1 2 n958-3 n691-2
0 n639 6 2 2 n649 n650
0 n680 6 2 2 n688 n689
0 n740 6 2 2 n748 n749
0 n778 6 2 2 n786 n787
0 n816 6 2 2 n824 n825
0 n882 6 2 2 n890 n891
0 n948 6 2 2 n956 n957
0 n995 6 2 2 n1003 n1004
2 n639-1 1 n639 
2 n639-2 1 n639 
2 n680-1 1 n680 
2 n680-2 1 n680 
2 n740-1 1 n740 
2 n740-2 1 n740 
2 n778-1 1 n778 
2 n778-2 1 n778 
2 n816-1 1 n816 
2 n816-2 1 n816 
2 n882-1 1 n882 
2 n882-2 1 n882 
2 n948-1 1 n948 
2 n948-2 1 n948 
2 n995-1 1 n995 
2 n995-2 1 n995 
0 n637 4 1 2 n638 n639-1
0 n647 5 2 1 n639-2
0 n678 4 1 2 n679 n680-1
0 n686 5 2 1 n680-2
0 n738 4 1 2 n739 n740-1
0 n746 5 2 1 n740-2
0 n776 4 1 2 n777 n778-1
0 n784 5 2 1 n778-2
0 n814 4 1 2 n815 n816-1
0 n822 5 2 1 n816-2
0 n880 4 1 2 n881 n882-1
0 n888 5 2 1 n882-2
0 n946 4 1 2 n947 n948-1
0 n954 5 2 1 n948-2
0 n993 4 1 2 n994 n995-1
0 n1001 5 2 1 n995-2
2 n647-1 1 n647 
2 n647-2 1 n647 
2 n686-1 1 n686 
2 n686-2 1 n686 
2 n746-1 1 n746 
2 n746-2 1 n746 
2 n784-1 1 n784 
2 n784-2 1 n784 
2 n822-1 1 n822 
2 n822-2 1 n822 
2 n888-1 1 n888 
2 n888-2 1 n888 
2 n954-1 1 n954 
2 n954-2 1 n954 
2 n1001-1 1 n1001 
2 n1001-2 1 n1001 
0 n646 4 1 2 n640-2 n647-1
0 n645 6 1 2 n648 n647-2
0 n685 4 1 2 n686-1 n641-2
0 n684 6 1 2 n687 n686-2
0 n745 4 1 2 n746-1 n641-3
0 n744 6 1 2 n747 n746-2
0 n783 4 1 2 n784-1 n641-4
0 n782 6 1 2 n785 n784-2
0 n821 4 1 2 n822-1 n641-5
0 n820 6 1 2 n823 n822-2
0 n887 4 1 2 n888-1 n641-6
0 n886 6 1 2 n889 n888-2
0 n953 4 1 2 n954-1 n641-7
0 n952 6 1 2 n955 n954-2
0 n1000 4 1 2 n641-8 n1001-1
0 n999 6 1 2 n1002 n1001-2
0 n642 6 2 2 n646 N233-1
0 n681 6 2 2 n685 N230-2
0 n741 6 2 2 n745 N228-2
0 n779 6 2 2 n783 N227-2
0 n817 6 2 2 n821 N226-2
0 n883 6 2 2 n887 N225-2
0 n949 6 2 2 n953 N229-2
0 n996 6 2 2 n1000 N231-2
2 n642-1 1 n642 
2 n642-2 1 n642 
2 n681-1 1 n681 
2 n681-2 1 n681 
2 n741-1 1 n741 
2 n741-2 1 n741 
2 n779-1 1 n779 
2 n779-2 1 n779 
2 n817-1 1 n817 
2 n817-2 1 n817 
2 n883-1 1 n883 
2 n883-2 1 n883 
2 n949-1 1 n949 
2 n949-2 1 n949 
2 n996-1 1 n996 
2 n996-2 1 n996 
0 n636 5 1 1 n642-1
0 n644 6 1 2 n645 n642-2
0 n677 5 1 1 n681-1
0 n683 6 1 2 n684 n681-2
0 n737 5 1 1 n741-1
0 n743 6 1 2 n744 n741-2
0 n775 5 1 1 n779-1
0 n781 6 1 2 n782 n779-2
0 n813 5 1 1 n817-1
0 n819 6 1 2 n820 n817-2
0 n879 5 1 1 n883-1
0 n885 6 1 2 n886 n883-2
0 n945 5 1 1 n949-1
0 n951 6 1 2 n952 n949-2
0 n992 5 1 1 n996-1
0 n998 6 1 2 n999 n996-2
0 n632 4 1 2 n636 n637
0 n630 6 1 2 n643 n644
0 n673 4 1 2 n677 n678
0 n671 6 1 2 n682 n683
0 n733 4 1 2 n737 n738
0 n731 6 1 2 n742 n743
0 n771 4 1 2 n775 n776
0 n769 6 1 2 n780 n781
0 n809 4 1 2 n813 n814
0 n807 6 1 2 n818 n819
0 n875 4 1 2 n879 n880
0 n873 6 1 2 n884 n885
0 n941 4 1 2 n945 n946
0 n939 6 1 2 n950 n951
0 n988 4 1 2 n992 n993
0 n986 6 1 2 n997 n998
0 n631 6 1 2 n632 n633
0 n672 6 1 2 n673 n674
0 n732 6 1 2 n733 n734
0 n770 6 1 2 n771 n772
0 n808 6 1 2 n809 n810
0 n874 6 1 2 n875 n876
0 n940 6 1 2 n941 n942
0 n987 6 1 2 n988 n989
0 n599 6 3 2 n630 n631
0 n580 6 4 2 n671 n672
0 n505 6 5 2 n731 n732
0 n503 6 2 2 n769 n770
0 n506 6 2 2 n807 n808
0 n504 6 3 2 n873 n874
0 n581 6 4 2 n939 n940
0 n560 6 5 2 n986 n987
2 n599-1 1 n599 
2 n599-2 1 n599 
2 n599-3 1 n599 
2 n580-1 1 n580 
2 n580-2 1 n580 
2 n580-3 1 n580 
2 n580-4 1 n580 
2 n505-1 1 n505 
2 n505-2 1 n505 
2 n505-3 1 n505 
2 n505-4 1 n505 
2 n505-5 1 n505 
2 n503-1 1 n503 
2 n503-2 1 n503 
2 n506-1 1 n506 
2 n506-2 1 n506 
2 n504-1 1 n504 
2 n504-2 1 n504 
2 n504-3 1 n504 
2 n581-1 1 n581 
2 n581-2 1 n581 
2 n581-3 1 n581 
2 n581-4 1 n581 
2 n560-1 1 n560 
2 n560-2 1 n560 
2 n560-3 1 n560 
2 n560-4 1 n560 
2 n560-5 1 n560 
0 n502 6 1 2 n503-1 n504-1
0 n499 4 1 2 n505-1 n506-1
0 n498 5 6 1 n581-1
0 n598 6 1 2 n599-1 n581-2
0 n595 4 1 2 n580-2 n560-3
0 n486 5 6 1 n599-2
0 n490 5 5 1 n560-4
0 n494 5 6 1 n580-3
0 n556 5 5 1 n505-3
0 n564 6 2 2 n599-3 n580-4
0 n555 5 7 1 n503-2
0 n522 5 8 1 n506-2
0 n539 5 7 1 n504-3
0 n628 4 1 2 n581-4 n560-5
2 n498-1 1 n498 
2 n498-2 1 n498 
2 n498-3 1 n498 
2 n498-4 1 n498 
2 n498-5 1 n498 
2 n498-6 1 n498 
2 n486-1 1 n486 
2 n486-2 1 n486 
2 n486-3 1 n486 
2 n486-4 1 n486 
2 n486-5 1 n486 
2 n486-6 1 n486 
2 n490-1 1 n490 
2 n490-2 1 n490 
2 n490-3 1 n490 
2 n490-4 1 n490 
2 n490-5 1 n490 
2 n494-1 1 n494 
2 n494-2 1 n494 
2 n494-3 1 n494 
2 n494-4 1 n494 
2 n494-5 1 n494 
2 n494-6 1 n494 
2 n556-1 1 n556 
2 n556-2 1 n556 
2 n556-3 1 n556 
2 n556-4 1 n556 
2 n556-5 1 n556 
2 n564-1 1 n564 
2 n564-2 1 n564 
2 n555-1 1 n555 
2 n555-2 1 n555 
2 n555-3 1 n555 
2 n555-4 1 n555 
2 n555-5 1 n555 
2 n555-6 1 n555 
2 n555-7 1 n555 
2 n522-1 1 n522 
2 n522-2 1 n522 
2 n522-3 1 n522 
2 n522-4 1 n522 
2 n522-5 1 n522 
2 n522-6 1 n522 
2 n522-7 1 n522 
2 n522-8 1 n522 
2 n539-1 1 n539 
2 n539-2 1 n539 
2 n539-3 1 n539 
2 n539-4 1 n539 
2 n539-5 1 n539 
2 n539-6 1 n539 
2 n539-7 1 n539 
0 n520 6 1 2 n522-1 n504-2
0 n562 6 1 2 n486-5 n494-5
0 n559 5 2 1 n564-1
0 n578 4 1 2 n498-6 n580-1
0 n613 4 1 2 n494-6 n581-3
0 n729 6 1 2 n555-6 n522-7
0 n538 4 3 2 n555-7 n522-8
2 n559-1 1 n559 
2 n559-2 1 n559 
2 n538-1 1 n538 
2 n538-2 1 n538 
2 n538-3 1 n538 
0 n536 7 1 2 n538-1 n539-1
0 n558 6 1 2 n559-1 n560-1
0 n563 4 1 2 n559-2 n560-2
0 n727 6 1 2 n505-4 n538-2
0 n730 4 1 2 n505-5 n538-3
0 n561 4 1 2 n563 n498-5
0 n728 4 1 2 n730 n539-7
0 n557 6 1 2 n561 n562
0 n726 6 1 2 n728 n729
0 n501 7 3 2 n557 n558
0 n597 7 3 2 n726 n727
2 n501-1 1 n501 
2 n501-2 1 n501 
2 n501-3 1 n501 
2 n597-1 1 n597 
2 n597-2 1 n597 
2 n597-3 1 n597 
0 n500 4 1 2 n502 n501-1
0 n537 4 1 2 n501-2 n505-2
0 n554 4 1 2 n501-3 n556-1
0 n596 4 1 2 n598 n597-1
0 n614 4 1 2 n490-5 n597-2
0 n629 4 1 2 n564-2 n597-3
0 n485 7 4 2 n499 n500
0 n526 7 4 2 n536 n537
0 n521 6 2 2 n554 n555-1
0 n585 7 4 2 n595 n596
0 n579 7 2 2 n614 n486-6
0 n618 7 4 2 n628 n629
2 n485-1 1 n485 
2 n485-2 1 n485 
2 n485-3 1 n485 
2 n485-4 1 n485 
2 n526-1 1 n526 
2 n526-2 1 n526 
2 n526-3 1 n526 
2 n526-4 1 n526 
2 n521-1 1 n521 
2 n521-2 1 n521 
2 n585-1 1 n585 
2 n585-2 1 n585 
2 n585-3 1 n585 
2 n585-4 1 n585 
2 n579-1 1 n579 
2 n579-2 1 n579 
2 n618-1 1 n618 
2 n618-2 1 n618 
2 n618-3 1 n618 
2 n618-4 1 n618 
0 n484 6 2 2 n485-1 n486-1
0 n489 6 2 2 n485-2 n490-1
0 n493 6 2 2 n485-3 n494-1
0 n497 6 2 2 n485-4 n498-1
0 n510 4 4 2 n520 n521-1
0 n525 6 2 2 n526-1 n486-3
0 n529 6 2 2 n526-2 n490-3
0 n532 6 2 2 n526-3 n494-3
0 n535 6 2 2 n526-4 n498-3
0 n553 4 1 2 n521-2 n522-2
0 n568 7 4 2 n578 n579-1
0 n584 6 2 2 n585-1 n556-3
0 n588 6 2 2 n585-2 n555-3
0 n591 6 2 2 n585-3 n522-4
0 n594 6 2 2 n585-4 n539-4
0 n603 7 4 2 n613 n579-2
0 n617 6 2 2 n556-5 n618-1
0 n621 6 2 2 n618-2 n555-5
0 n624 6 2 2 n618-3 n522-6
0 n627 6 2 2 n618-4 n539-6
0 n543 7 4 2 n553 n539-2
2 n484-1 1 n484 
2 n484-2 1 n484 
2 n489-1 1 n489 
2 n489-2 1 n489 
2 n493-1 1 n493 
2 n493-2 1 n493 
2 n497-1 1 n497 
2 n497-2 1 n497 
2 n510-1 1 n510 
2 n510-2 1 n510 
2 n510-3 1 n510 
2 n510-4 1 n510 
2 n525-1 1 n525 
2 n525-2 1 n525 
2 n529-1 1 n529 
2 n529-2 1 n529 
2 n532-1 1 n532 
2 n532-2 1 n532 
2 n535-1 1 n535 
2 n535-2 1 n535 
2 n568-1 1 n568 
2 n568-2 1 n568 
2 n568-3 1 n568 
2 n568-4 1 n568 
2 n584-1 1 n584 
2 n584-2 1 n584 
2 n588-1 1 n588 
2 n588-2 1 n588 
2 n591-1 1 n591 
2 n591-2 1 n591 
2 n594-1 1 n594 
2 n594-2 1 n594 
2 n603-1 1 n603 
2 n603-2 1 n603 
2 n603-3 1 n603 
2 n603-4 1 n603 
2 n617-1 1 n617 
2 n617-2 1 n617 
2 n621-1 1 n621 
2 n621-2 1 n621 
2 n624-1 1 n624 
2 n624-2 1 n624 
2 n627-1 1 n627 
2 n627-2 1 n627 
0 n483 6 1 2 N218-1 n484-1
0 n482 3 1 2 N218-2 n484-2
0 n488 6 1 2 N211-1 n489-1
0 n487 3 1 2 N211-2 n489-2
0 n492 6 1 2 N204-1 n493-1
0 n491 3 1 2 N204-2 n493-2
0 n496 6 1 2 N197-1 n497-1
0 n495 3 1 2 N197-2 n497-2
0 n509 6 2 2 n510-1 n486-2
0 n513 6 2 2 n510-2 n490-2
0 n516 6 2 2 n510-3 n494-2
0 n519 6 2 2 n510-4 n498-2
0 n524 6 1 2 N162-1 n525-1
0 n523 3 1 2 N162-2 n525-2
0 n528 6 1 2 N155-1 n529-1
0 n527 3 1 2 N155-2 n529-2
0 n531 6 1 2 N148-1 n532-1
0 n530 3 1 2 N148-2 n532-2
0 n534 6 1 2 N141-1 n535-1
0 n533 3 1 2 N141-2 n535-2
0 n567 6 2 2 n568-1 n556-2
0 n571 6 2 2 n568-2 n555-2
0 n574 6 2 2 n568-3 n522-3
0 n577 6 2 2 n568-4 n539-3
0 n583 6 1 2 N78-1 n584-1
0 n582 3 1 2 N78-2 n584-2
0 n587 6 1 2 N71-1 n588-1
0 n586 3 1 2 N71-2 n588-2
0 n590 6 1 2 N64-1 n591-1
0 n589 3 1 2 N64-2 n591-2
0 n593 6 1 2 N57-1 n594-1
0 n592 3 1 2 N57-2 n594-2
0 n602 6 2 2 n603-1 n556-4
0 n606 6 2 2 n603-2 n555-4
0 n609 6 2 2 n603-3 n522-5
0 n612 6 2 2 n603-4 n539-5
0 n616 6 1 2 N22-1 n617-1
0 n615 3 1 2 N22-2 n617-2
0 n620 6 1 2 N15-1 n621-1
0 n619 3 1 2 N15-2 n621-2
0 n623 6 1 2 N8-1 n624-1
0 n622 3 1 2 N8-2 n624-2
0 n626 6 1 2 N1-1 n627-1
0 n625 3 1 2 N1-2 n627-2
2 n543-1 1 n543 
2 n543-2 1 n543 
2 n543-3 1 n543 
2 n543-4 1 n543 
3 N1355 6 0 2 n482 n483
3 N1354 6 0 2 n487 n488
3 N1353 6 0 2 n491 n492
3 N1352 6 0 2 n495 n496
3 N1347 6 0 2 n523 n524
3 N1346 6 0 2 n527 n528
3 N1345 6 0 2 n530 n531
3 N1344 6 0 2 n533 n534
0 n542 6 2 2 n543-1 n486-4
0 n546 6 2 2 n543-2 n490-4
0 n549 6 2 2 n543-3 n494-4
0 n552 6 2 2 n543-4 n498-4
3 N1335 6 0 2 n582 n583
3 N1334 6 0 2 n586 n587
3 N1333 6 0 2 n589 n590
3 N1332 6 0 2 n592 n593
3 N1327 6 0 2 n615 n616
3 N1326 6 0 2 n619 n620
3 N1325 6 0 2 n622 n623
3 N1324 6 0 2 n625 n626
2 n509-1 1 n509 
2 n509-2 1 n509 
2 n513-1 1 n513 
2 n513-2 1 n513 
2 n516-1 1 n516 
2 n516-2 1 n516 
2 n519-1 1 n519 
2 n519-2 1 n519 
2 n567-1 1 n567 
2 n567-2 1 n567 
2 n571-1 1 n571 
2 n571-2 1 n571 
2 n574-1 1 n574 
2 n574-2 1 n574 
2 n577-1 1 n577 
2 n577-2 1 n577 
2 n602-1 1 n602 
2 n602-2 1 n602 
2 n606-1 1 n606 
2 n606-2 1 n606 
2 n609-1 1 n609 
2 n609-2 1 n609 
2 n612-1 1 n612 
2 n612-2 1 n612 
0 n508 6 1 2 N190-1 n509-1
0 n507 3 1 2 N190-2 n509-2
0 n512 6 1 2 N183-1 n513-1
0 n511 3 1 2 N183-2 n513-2
0 n515 6 1 2 N176-1 n516-1
0 n514 3 1 2 N176-2 n516-2
0 n518 6 1 2 N169-1 n519-1
0 n517 3 1 2 N169-2 n519-2
0 n566 6 1 2 N106-1 n567-1
0 n565 3 1 2 N106-2 n567-2
0 n570 6 1 2 N99-1 n571-1
0 n569 3 1 2 N99-2 n571-2
0 n573 6 1 2 N92-1 n574-1
0 n572 3 1 2 N92-2 n574-2
0 n576 6 1 2 N85-1 n577-1
0 n575 3 1 2 N85-2 n577-2
0 n601 6 1 2 N50-1 n602-1
0 n600 3 1 2 N50-2 n602-2
0 n605 6 1 2 N43-1 n606-1
0 n604 3 1 2 N43-2 n606-2
0 n608 6 1 2 N36-1 n609-1
0 n607 3 1 2 N36-2 n609-2
0 n611 6 1 2 N29-1 n612-1
0 n610 3 1 2 N29-2 n612-2
2 n542-1 1 n542 
2 n542-2 1 n542 
2 n546-1 1 n546 
2 n546-2 1 n546 
2 n549-1 1 n549 
2 n549-2 1 n549 
2 n552-1 1 n552 
2 n552-2 1 n552 
3 N1351 6 0 2 n507 n508
3 N1350 6 0 2 n511 n512
3 N1349 6 0 2 n514 n515
3 N1348 6 0 2 n517 n518
0 n541 6 1 2 N134-1 n542-1
0 n540 3 1 2 N134-2 n542-2
0 n545 6 1 2 N127-1 n546-1
0 n544 3 1 2 N127-2 n546-2
0 n548 6 1 2 N120-1 n549-1
0 n547 3 1 2 N120-2 n549-2
0 n551 6 1 2 N113-1 n552-1
0 n550 3 1 2 N113-2 n552-2
3 N1339 6 0 2 n565 n566
3 N1338 6 0 2 n569 n570
3 N1337 6 0 2 n572 n573
3 N1336 6 0 2 n575 n576
3 N1331 6 0 2 n600 n601
3 N1330 6 0 2 n604 n605
3 N1329 6 0 2 n607 n608
3 N1328 6 0 2 n610 n611
3 N1343 6 0 2 n540 n541
3 N1342 6 0 2 n544 n545
3 N1341 6 0 2 n547 n548
3 N1340 6 0 2 n550 n551
