1 1 0 1 0 
1 2 0 1 0 
1 3 0 1 0 
1 4 0 1 0 
1 5 0 1 0 
0 6 7 2 1 1 
2 7 1 6 
2 8 1 6 
0 9 7 2 1 2 
2 10 1 9 
2 11 1 9 
0 12 7 2 1 3 
2 13 1 12 
2 14 1 12 
0 15 7 2 1 4 
2 16 1 15 
2 17 1 15 
0 18 7 2 1 5 
2 19 1 18 
2 20 1 18 
0 21 5 1 1 7 
0 22 3 1 2 10 13 
0 23 6 2 2 11 14 
2 24 1 23 
2 25 1 23 
0 26 6 2 2 22 24 
2 27 1 26 
2 28 1 26 
0 29 6 1 2 21 27 
0 30 5 1 1 28 
0 31 6 2 2 8 30 
2 32 1 31 
2 33 1 31 
0 34 6 2 2 33 25 
2 35 1 34 
2 36 1 34 
0 37 5 1 1 35 
0 38 3 1 2 16 19 
0 39 6 2 2 17 20 
2 40 1 39 
2 41 1 39 
0 42 6 2 2 38 40 
2 43 1 42 
2 44 1 42 
0 45 6 1 2 37 43 
0 46 5 1 1 44 
0 47 6 2 2 36 46 
2 48 1 47 
2 49 1 47 
3 50 7 0 2 29 32 
3 51 7 0 2 45 48 
3 52 6 0 2 49 41 
