1 1 0 2 0 
2 2 1 1  
2 3 1 1  
1 4 0 3 0 
2 5 1 4  
2 6 1 4  
2 7 1 4  
1 8 0 2 0 
2 9 1 8  
2 10 1 8  
1 11 0 2 0 
2 12 1 11  
2 13 1 11  
1 14 0 2 0 
2 15 1 14  
2 16 1 14  
1 17 0 3 0 
2 18 1 17  
2 19 1 17  
2 20 1 17  
1 21 0 2 0 
2 22 1 21  
2 23 1 21  
1 24 0 2 0 
2 25 1 24  
2 26 1 24  
1 27 0 2 0 
2 28 1 27  
2 29 1 27  
1 30 0 3 0 
2 31 1 30  
2 32 1 30  
2 33 1 30  
1 34 0 2 0 
2 35 1 34  
2 36 1 34  
1 37 0 2 0 
2 38 1 37  
2 39 1 37  
1 40 0 2 0 
2 41 1 40  
2 42 1 40  
1 43 0 3 0 
2 44 1 43  
2 45 1 43  
2 46 1 43  
1 47 0 2 0 
2 48 1 47  
2 49 1 47  
1 50 0 2 0 
2 51 1 50  
2 52 1 50  
1 53 0 2 0 
2 54 1 53  
2 55 1 53  
1 56 0 3 0 
2 57 1 56  
2 58 1 56  
2 59 1 56  
1 60 0 2 0 
2 61 1 60  
2 62 1 60  
1 63 0 2 0 
2 64 1 63  
2 65 1 63  
1 66 0 2 0 
2 67 1 66  
2 68 1 66  
1 69 0 3 0 
2 70 1 69  
2 71 1 69  
2 72 1 69  
1 73 0 2 0 
2 74 1 73  
2 75 1 73  
1 76 0 2 0 
2 77 1 76  
2 78 1 76  
1 79 0 2 0 
2 80 1 79  
2 81 1 79  
1 82 0 3 0 
2 83 1 82  
2 84 1 82  
2 85 1 82  
1 86 0 2 0 
2 87 1 86  
2 88 1 86  
1 89 0 2 0 
2 90 1 89  
2 91 1 89  
1 92 0 2 0 
2 93 1 92  
2 94 1 92  
1 95 0 3 0 
2 96 1 95  
2 97 1 95  
2 98 1 95  
1 99 0 2 0 
2 100 1 99  
2 101 1 99  
1 102 0 2 0 
2 103 1 102  
2 104 1 102  
1 105 0 2 0 
2 106 1 105  
2 107 1 105  
1 108 0 3 0 
2 109 1 108  
2 110 1 108  
2 111 1 108  
1 112 0 2 0 
2 113 1 112  
2 114 1 112  
1 115 0 2 0 
2 116 1 115  
2 117 1 115  
0 118 5 1 1 2 
0 119 5 2 1 5 
2 120 1 119  
2 121 1 119  
0 122 5 1 1 12 
0 123 5 2 1 18 
2 124 1 123  
2 125 1 123  
0 126 5 1 1 25 
0 127 5 2 1 31 
2 128 1 127  
2 129 1 127  
0 130 5 1 1 38 
0 131 5 2 1 44 
2 132 1 131  
2 133 1 131  
0 134 5 1 1 51 
0 135 5 2 1 57 
2 136 1 135  
2 137 1 135  
0 138 5 1 1 64 
0 139 5 2 1 70 
2 140 1 139  
2 141 1 139  
0 142 5 1 1 77 
0 143 5 2 1 83 
2 144 1 143  
2 145 1 143  
0 146 5 1 1 90 
0 147 5 2 1 96 
2 148 1 147  
2 149 1 147  
0 150 5 1 1 103 
0 151 5 2 1 109 
2 152 1 151  
2 153 1 151  
0 154 6 2 2 118 6 
2 155 1 154  
2 156 1 154  
0 157 4 1 2 9 120 
0 158 4 1 2 15 121 
0 159 6 2 2 122 19 
2 160 1 159  
2 161 1 159  
0 162 6 2 2 126 32 
2 163 1 162  
2 164 1 162  
0 165 6 2 2 130 45 
2 166 1 165  
2 167 1 165  
0 168 6 2 2 134 58 
2 169 1 168  
2 170 1 168  
0 171 6 2 2 138 71 
2 172 1 171  
2 173 1 171  
0 174 6 2 2 142 84 
2 175 1 174  
2 176 1 174  
0 177 6 2 2 146 97 
2 178 1 177  
2 179 1 177  
0 180 6 2 2 150 110 
2 181 1 180  
2 182 1 180  
0 183 4 1 2 22 124 
0 184 4 1 2 28 125 
0 185 4 1 2 35 128 
0 186 4 1 2 41 129 
0 187 4 1 2 48 132 
0 188 4 1 2 54 133 
0 189 4 1 2 61 136 
0 190 4 1 2 67 137 
0 191 4 1 2 74 140 
0 192 4 1 2 80 141 
0 193 4 1 2 87 144 
0 194 4 1 2 93 145 
0 195 4 1 2 100 148 
0 196 4 1 2 106 149 
0 197 4 1 2 113 152 
0 198 4 1 2 116 153 
0 199 7 3 9 155 160 163 166 169 172 175 178 181 
2 200 1 199  
2 201 1 199  
2 202 1 199  
0 203 5 9 1 200 
2 204 1 203  
2 205 1 203  
2 206 1 203  
2 207 1 203  
2 208 1 203  
2 209 1 203  
2 210 1 203  
2 211 1 203  
2 212 1 203  
0 213 5 9 1 201 
2 214 1 213  
2 215 1 213  
2 216 1 213  
2 217 1 213  
2 218 1 213  
2 219 1 213  
2 220 1 213  
2 221 1 213  
2 222 1 213  
3 223 5 0 1 202 
0 224 2 2 2 204 156 
2 225 1 224  
2 226 1 224  
0 227 2 2 2 205 161 
2 228 1 227  
2 229 1 227  
0 230 2 2 2 206 164 
2 231 1 230  
2 232 1 230  
0 233 2 2 2 207 167 
2 234 1 233  
2 235 1 233  
0 236 2 2 2 208 170 
2 237 1 236  
2 238 1 236  
0 239 2 2 2 209 173 
2 240 1 239  
2 241 1 239  
0 242 6 1 2 3 214 
0 243 2 2 2 210 176 
2 244 1 243  
2 245 1 243  
0 246 6 1 2 215 13 
0 247 2 2 2 211 179 
2 248 1 247  
2 249 1 247  
0 250 6 1 2 216 26 
0 251 2 2 2 212 182 
2 252 1 251  
2 253 1 251  
0 254 6 1 2 217 39 
0 255 6 1 2 218 52 
0 256 6 1 2 219 65 
0 257 6 1 2 220 78 
0 258 6 1 2 221 91 
0 259 6 1 2 222 104 
0 260 6 2 2 225 157 
2 261 1 260  
2 262 1 260  
0 263 6 1 2 226 158 
0 264 6 2 2 228 183 
2 265 1 264  
2 266 1 264  
0 267 6 2 2 231 185 
2 268 1 267  
2 269 1 267  
0 270 6 2 2 234 187 
2 271 1 270  
2 272 1 270  
0 273 6 2 2 237 189 
2 274 1 273  
2 275 1 273  
0 276 6 2 2 240 191 
2 277 1 276  
2 278 1 276  
0 279 6 2 2 244 193 
2 280 1 279  
2 281 1 279  
0 282 6 2 2 248 195 
2 283 1 282  
2 284 1 282  
0 285 6 2 2 252 197 
2 286 1 285  
2 287 1 285  
0 288 6 1 2 229 184 
0 289 6 1 2 232 186 
0 290 6 1 2 235 188 
0 291 6 1 2 238 190 
0 292 6 1 2 241 192 
0 293 6 1 2 245 194 
0 294 6 1 2 249 196 
0 295 6 1 2 253 198 
0 296 7 3 9 261 265 268 271 274 277 280 283 286 
2 297 1 296  
2 298 1 296  
2 299 1 296  
0 300 5 1 1 263 
0 301 5 1 1 288 
0 302 5 1 1 289 
0 303 5 1 1 290 
0 304 5 1 1 291 
0 305 5 1 1 292 
0 306 5 1 1 293 
0 307 5 1 1 294 
0 308 5 1 1 295 
0 309 5 9 1 297 
2 310 1 309  
2 311 1 309  
2 312 1 309  
2 313 1 309  
2 314 1 309  
2 315 1 309  
2 316 1 309  
2 317 1 309  
2 318 1 309  
0 319 5 9 1 298 
2 320 1 319  
2 321 1 319  
2 322 1 319  
2 323 1 319  
2 324 1 319  
2 325 1 319  
2 326 1 319  
2 327 1 319  
2 328 1 319  
3 329 5 0 1 299 
0 330 2 1 2 310 262 
0 331 2 1 2 311 266 
0 332 2 1 2 312 269 
0 333 2 1 2 313 272 
0 334 6 1 2 10 320 
0 335 2 1 2 314 275 
0 336 6 1 2 321 23 
0 337 2 1 2 315 278 
0 338 6 1 2 322 36 
0 339 2 1 2 316 281 
0 340 6 1 2 323 49 
0 341 2 1 2 317 284 
0 342 6 1 2 324 62 
0 343 2 1 2 318 287 
0 344 6 1 2 325 75 
0 345 6 1 2 326 88 
0 346 6 1 2 327 101 
0 347 6 1 2 328 114 
0 348 6 1 2 330 300 
0 349 6 1 2 331 301 
0 350 6 1 2 332 302 
0 351 6 1 2 333 303 
0 352 6 1 2 335 304 
0 353 6 1 2 337 305 
0 354 6 1 2 339 306 
0 355 6 1 2 341 307 
0 356 6 1 2 343 308 
0 357 7 2 9 348 349 350 351 352 353 354 355 356 
2 358 1 357  
2 359 1 357  
0 360 5 9 1 358 
2 361 1 360  
2 362 1 360  
2 363 1 360  
2 364 1 360  
2 365 1 360  
2 366 1 360  
2 367 1 360  
2 368 1 360  
2 369 1 360  
3 370 5 0 1 359 
0 371 6 1 2 16 361 
0 372 6 1 2 362 29 
0 373 6 1 2 363 42 
0 374 6 1 2 364 55 
0 375 6 1 2 365 68 
0 376 6 1 2 366 81 
0 377 6 1 2 367 94 
0 378 6 1 2 368 107 
0 379 6 1 2 369 117 
0 380 6 1 4 7 242 334 371 
0 381 6 4 4 246 336 372 20 
2 382 1 381  
2 383 1 381  
2 384 1 381  
2 385 1 381  
0 386 6 6 4 250 338 373 33 
2 387 1 386  
2 388 1 386  
2 389 1 386  
2 390 1 386  
2 391 1 386  
2 392 1 386  
0 393 6 5 4 254 340 374 46 
2 394 1 393  
2 395 1 393  
2 396 1 393  
2 397 1 393  
2 398 1 393  
0 399 6 4 4 255 342 375 59 
2 400 1 399  
2 401 1 399  
2 402 1 399  
2 403 1 399  
0 404 6 2 4 256 344 376 72 
2 405 1 404  
2 406 1 404  
0 407 6 3 4 257 345 377 85 
2 408 1 407  
2 409 1 407  
2 410 1 407  
0 411 6 2 4 258 346 378 98 
2 412 1 411  
2 413 1 411  
0 414 6 1 4 259 347 379 111 
0 415 5 1 1 380 
0 416 7 1 8 382 387 394 400 405 408 412 414 
0 417 5 1 1 395 
0 418 5 1 1 406 
0 419 5 1 1 409 
0 420 5 1 1 413 
3 421 4 0 2 415 416 
0 422 6 2 2 388 417 
2 423 1 422  
2 424 1 422  
0 425 6 2 4 389 396 418 401 
2 426 1 425  
2 427 1 425  
0 428 6 1 3 402 397 419 
0 429 6 1 4 390 398 410 420 
3 430 6 0 4 383 391 423 403 
3 431 6 0 4 384 392 426 428 
3 432 6 0 4 385 424 427 429 
