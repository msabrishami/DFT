1 1 0 11 0
1 13 0 6 0
1 20 0 12 0
1 33 0 7 0
1 41 0 3 0
1 45 0 4 0
1 50 0 7 0
1 58 0 9 0
1 68 0 8 0
1 77 0 9 0
1 87 0 9 0
1 97 0 9 0
1 107 0 8 0
1 116 0 7 0
1 124 0 1 0
1 125 0 2 0
1 128 0 3 0
1 132 0 4 0
1 137 0 5 0
1 143 0 6 0
1 150 0 8 0
1 159 0 9 0
1 169 0 9 0
1 179 0 10 0
1 190 0 9 0
1 200 0 12 0
1 213 0 8 0
1 222 0 1 0
1 223 0 2 0
1 226 0 5 0
1 232 0 5 0
1 238 0 5 0
1 244 0 5 0
1 250 0 6 0
1 257 0 6 0
1 264 0 5 0
1 270 0 3 0
1 274 0 8 0
1 283 0 10 0
1 294 0 8 0
1 303 0 7 0
1 311 0 5 0
1 317 0 4 0
1 322 0 3 0
1 326 0 2 0
1 329 0 1 0
1 330 0 12 0
1 343 0 5 0
1 349 0 1 0
1 350 0 2 0
0 655 9 9 1 51
0 665 5 4 1 52
0 670 9 8 1 59
0 679 5 3 1 60
0 683 9 2 1 69
0 686 5 3 1 70
0 690 9 8 1 71
0 699 9 2 1 78
0 702 5 3 1 79
0 706 9 8 1 80
0 715 9 8 1 88
0 724 5 2 1 89
0 727 9 8 1 98
0 736 5 3 1 99
0 740 9 8 1 108
0 749 5 3 1 109
0 753 9 9 1 117
0 763 5 4 1 118
0 768 3 1 2 258 265
0 769 5 2 1 2
0 772 9 6 1 3
0 779 5 2 1 4
0 782 9 3 1 14
0 786 5 6 1 15
0 793 7 1 2 16 21
0 794 5 3 1 22
0 798 9 4 1 23
0 803 5 16 1 24
0 820 5 1 1 34
0 821 9 3 1 35
0 825 5 3 1 36
0 829 7 2 2 37 42
0 832 5 2 1 43
0 835 3 1 2 44 46
0 836 9 2 1 47
0 839 5 2 1 48
0 842 5 2 1 53
0 845 9 2 1 61
0 848 5 2 1 62
0 851 9 2 1 72
0 854 5 3 1 73
0 858 9 2 1 90
0 861 5 2 1 91
0 864 9 2 1 100
0 867 5 2 1 101
0 870 5 3 1 110
0 874 9 2 1 5
0 877 9 2 1 74
0 880 9 2 1 111
0 883 5 2 1 25
0 886 9 2 1 191
0 889 5 1 1 201
0 890 7 1 2 26 202
0 891 6 1 2 27 203
0 892 7 2 2 28 180
0 895 5 1 1 29
0 896 3 16 2 349 38
0 913 6 1 2 6 17
0 914 6 1 3 7 30 39
0 915 5 1 1 31
0 916 5 1 1 40
0 917 9 2 1 181
0 920 5 2 1 214
0 923 9 2 1 344
0 926 9 2 1 227
0 929 9 2 1 233
0 932 9 2 1 239
0 935 9 2 1 245
0 938 9 2 1 251
0 941 9 2 1 259
0 944 9 2 1 266
0 947 9 2 1 271
0 950 9 2 1 54
0 953 9 2 1 63
0 956 9 2 1 64
0 959 9 2 1 102
0 962 9 2 1 103
0 965 9 2 1 331
0 1067 7 1 2 252 768
0 1117 3 16 2 820 32
0 1179 3 1 2 895 170
0 1196 5 1 1 793
0 1197 3 4 2 915 8
0 1202 7 16 2 913 914
0 1219 3 4 2 916 9
0 1250 7 1 3 504 508 512
0 1251 6 1 2 228 353
0 1252 6 1 2 234 366
0 1253 6 1 2 240 382
0 1254 6 1 2 246 395
0 1255 6 1 2 253 403
0 1256 6 1 2 260 413
0 1257 6 1 2 267 424
0 1258 6 1 2 272 435
0 1259 5 1 1 560
0 1260 5 1 1 562
0 1261 5 1 1 564
0 1262 5 1 1 566
0 1263 6 1 2 374 379
0 1264 6 2 2 421 432
0 1267 6 1 2 377 390
0 1268 9 2 1 362
0 1271 5 1 1 578
0 1272 5 1 1 582
0 1273 9 2 1 502
0 1276 9 2 1 503
0 1279 9 2 1 458
0 1298 9 3 1 493
0 1302 9 3 1 498
0 1306 7 8 2 456 835
0 1315 7 6 3 457 500 499
0 1322 7 2 2 448 501
0 1325 7 2 3 450 461 470
0 1328 6 2 3 451 462 471
0 1331 6 2 2 452 463
0 1334 9 2 1 526
0 1337 6 1 3 459 467 49
0 1338 6 1 3 505 509 513
0 1339 5 1 1 580
0 1340 7 2 3 517 521 523
0 1343 6 1 3 518 522 524
0 1344 5 1 1 584
0 1345 5 1 1 474
0 1346 5 1 1 475
0 1347 5 1 1 476
0 1348 5 1 1 477
0 1349 5 1 1 478
0 1350 5 1 1 479
0 1351 5 1 1 480
0 1352 5 1 1 481
0 1353 3 4 2 532 534
0 1358 4 4 2 533 535
0 1363 9 2 1 536
0 1366 5 2 1 537
0 1369 9 14 1 490
0 1384 9 16 1 494
0 1401 5 1 1 538
0 1402 5 1 1 539
0 1403 5 1 1 540
0 1404 5 1 1 541
0 1405 5 1 1 542
0 1406 5 1 1 543
0 1407 5 1 1 544
0 1408 5 1 1 545
0 1409 3 16 2 10 1196
0 1426 5 1 1 496
0 1427 5 1 1 497
0 1452 7 6 3 449 460 468
0 1459 5 1 1 554
0 1460 5 1 1 586
0 1461 3 2 2 556 558
0 1464 4 2 2 557 559
0 1467 5 1 1 568
0 1468 5 1 1 570
0 1469 5 1 1 572
0 1470 5 1 1 574
0 1471 9 2 1 375
0 1474 5 1 1 576
0 1475 9 2 1 380
0 1478 9 2 1 392
0 1481 9 2 1 411
0 1484 9 2 1 422
0 1487 9 2 1 433
0 1490 9 2 1 444
0 1493 9 2 1 528
0 1496 9 2 1 529
0 1499 9 2 1 530
0 1502 9 2 1 531
0 1505 6 1 2 393 1250
0 1507 7 1 4 1251 1252 1253 1254
0 1508 7 1 4 1255 1256 1257 1258
0 1509 6 1 2 563 1259
0 1510 6 1 2 561 1260
0 1511 6 1 2 567 1261
0 1512 6 1 2 565 1262
0 1520 7 3 2 354 1263
0 1562 7 16 2 527 1337
0 1579 5 1 1 588
0 1580 7 1 2 482 589
0 1581 7 1 2 1338 1345
0 1582 5 1 1 590
0 1583 7 1 2 483 591
0 1584 5 1 1 592
0 1585 7 1 2 484 593
0 1586 7 1 2 514 1347
0 1587 5 1 1 594
0 1588 7 1 2 485 595
0 1589 7 1 2 81 1348
0 1590 5 1 1 596
0 1591 7 1 2 486 597
0 1592 7 1 2 1343 1349
0 1593 5 1 1 598
0 1594 7 1 2 487 599
0 1595 5 1 1 600
0 1596 7 1 2 488 601
0 1597 7 1 2 525 1351
0 1598 5 1 1 602
0 1599 7 1 2 489 603
0 1600 7 1 2 119 1352
0 1643 7 1 2 222 1401
0 1644 7 1 2 224 1402
0 1645 7 1 2 229 1403
0 1646 7 1 2 235 1404
0 1647 7 1 2 241 1405
0 1648 7 1 2 247 1406
0 1649 7 1 2 254 1407
0 1650 7 1 2 261 1408
0 1667 7 2 3 11 18 1426
0 1670 7 2 3 12 19 1427
0 1673 5 1 1 608
0 1674 5 1 1 609
0 1675 5 1 1 610
0 1676 5 1 1 611
0 1677 5 1 1 612
0 1678 5 1 1 613
0 1679 5 1 1 614
0 1680 5 1 1 615
0 1691 6 1 2 571 1467
0 1692 6 1 2 569 1468
0 1693 6 1 2 575 1469
0 1694 6 1 2 573 1470
3 1713 5 0 1 1505
0 1714 7 1 2 92 628
0 1715 6 2 2 1509 1510
0 1718 6 2 2 1511 1512
0 1721 6 1 2 1507 1508
0 1722 7 2 2 445 671
0 1725 6 1 2 446 672
0 1726 5 1 1 630
0 1727 6 1 2 773 1271
0 1728 5 1 1 774
0 1729 7 1 2 378 631
0 1730 6 1 2 777 1272
0 1731 5 1 1 778
0 1735 6 1 2 93 629
0 1736 5 1 1 632
0 1737 5 1 1 634
0 1738 6 8 2 661 491
0 1747 6 8 2 662 495
0 1756 6 4 3 453 636 472
0 1761 6 2 4 454 464 473 641
0 1764 6 1 2 775 1339
0 1765 5 1 1 776
0 1766 6 1 2 780 1344
0 1767 5 1 1 781
0 1768 5 1 1 663
0 1769 5 1 1 668
0 1770 5 1 1 666
0 1787 7 1 2 506 1579
0 1788 7 1 2 151 1580
0 1789 7 1 2 510 1582
0 1790 7 1 2 160 1583
0 1791 7 1 2 82 1584
0 1792 7 1 2 55 1585
0 1793 7 1 2 515 1587
0 1794 7 1 2 507 1588
0 1795 7 1 2 519 1590
0 1796 7 1 2 511 1591
0 1797 7 1 2 112 1593
0 1798 7 1 2 83 1594
0 1799 7 1 2 120 1595
0 1800 7 1 2 516 1596
0 1801 7 1 2 284 1598
0 1802 7 1 2 520 1599
0 1803 7 2 2 204 682
0 1806 7 2 2 889 684
0 1809 7 2 2 890 685
0 1812 7 2 2 891 687
0 1815 6 2 2 638 642
0 1818 6 2 2 492 643
0 1821 6 2 3 455 637 1179
0 1824 6 8 3 465 469 639
0 1833 6 8 2 466 640
0 1842 5 1 1 688
0 1843 5 1 1 689
0 1844 5 1 1 691
0 1845 5 1 1 692
0 1846 5 1 1 693
0 1847 5 1 1 694
0 1848 5 1 1 695
0 1849 5 1 1 705
0 1850 7 1 2 707 546
0 1851 5 1 1 708
0 1852 7 1 2 709 547
0 1853 5 1 1 710
0 1854 7 1 2 711 548
0 1855 5 1 1 712
0 1856 7 1 2 713 549
0 1857 5 1 1 714
0 1858 7 1 2 716 550
0 1859 5 1 1 717
0 1860 7 1 2 718 551
0 1861 5 1 1 719
0 1862 7 1 2 720 552
0 1863 5 1 1 721
0 1864 7 1 2 722 553
0 1869 7 1 2 616 723
0 1870 4 2 2 56 725
0 1873 5 1 1 644
0 1874 7 1 2 617 726
0 1875 4 2 2 65 728
0 1878 5 1 1 645
0 1879 7 1 2 618 729
0 1880 4 2 2 75 730
0 1883 5 1 1 646
0 1884 7 1 2 619 731
0 1885 4 2 2 84 732
0 1888 5 1 1 647
0 1889 7 1 2 620 733
0 1890 4 2 2 94 734
0 1893 5 1 1 659
0 1894 7 1 2 621 735
0 1895 4 2 2 104 737
0 1898 5 1 1 652
0 1899 7 1 2 622 738
0 1900 4 2 2 113 739
0 1903 5 1 1 653
0 1904 7 1 2 623 741
0 1905 4 2 2 121 742
0 1908 5 1 1 654
0 1909 7 2 2 743 215
0 1912 6 1 2 744 216
0 1913 7 3 3 745 217 345
0 1917 6 4 3 746 218 346
0 1922 7 3 3 747 219 347
0 1926 6 3 3 748 220 348
0 1930 9 2 1 752
0 1933 6 2 2 1691 1692
0 1936 6 2 2 1693 1694
0 1939 5 1 1 755
0 1940 6 1 2 756 1474
0 1941 5 1 1 757
0 1942 5 1 1 759
0 1943 5 1 1 761
0 1944 5 1 1 764
0 1945 5 1 1 766
0 1946 5 1 1 770
3 1947 5 0 1 1714
0 1960 6 1 2 579 1728
0 1961 6 1 2 583 1731
0 1966 7 1 2 783 635
0 1981 6 1 2 581 1765
0 1982 6 1 2 585 1767
0 1983 7 2 2 1067 1768
0 1986 3 1 3 1581 1787 1788
0 1987 3 1 3 1586 1791 1792
0 1988 3 1 3 1589 1793 1794
0 1989 3 1 3 1592 1795 1796
0 1990 3 1 3 1597 1799 1800
0 1991 3 1 3 1600 1801 1802
0 2022 7 1 2 85 1849
0 2023 7 1 2 225 1850
0 2024 7 1 2 95 1851
0 2025 7 1 2 230 1852
0 2026 7 1 2 105 1853
0 2027 7 1 2 236 1854
0 2028 7 1 2 114 1855
0 2029 7 1 2 242 1856
0 2030 7 1 2 122 1857
0 2031 7 1 2 248 1858
0 2032 7 1 2 285 1859
0 2033 7 1 2 255 1860
0 2034 7 1 2 295 1861
0 2035 7 1 2 262 1862
0 2036 7 1 2 304 1863
0 2037 7 1 2 268 1864
0 2038 9 4 1 807
0 2043 5 8 1 808
0 2052 9 4 1 809
0 2057 5 8 1 810
0 2068 7 2 3 57 604 1869
0 2073 7 2 3 66 605 1874
0 2078 7 2 3 76 606 1879
0 2083 7 2 3 86 607 1884
0 2088 7 2 3 96 624 1889
0 2093 7 2 3 106 625 1894
0 2098 7 2 3 115 626 1899
0 2103 7 2 3 123 627 1904
0 2121 5 1 1 787
0 2122 5 1 1 788
0 2123 5 1 1 789
0 2124 5 1 1 790
0 2125 5 1 1 791
0 2126 5 1 1 792
0 2127 5 1 1 795
0 2128 5 1 1 796
0 2133 6 1 2 577 1939
0 2134 6 1 2 760 1941
0 2135 6 1 2 758 1942
0 2136 6 1 2 765 1943
0 2137 6 1 2 762 1944
0 2138 6 1 2 771 1945
0 2139 6 1 2 767 1946
0 2141 5 1 1 945
0 2142 5 1 1 948
0 2143 5 1 1 817
0 2144 7 1 2 818 828
0 2145 5 1 1 830
0 2146 6 1 2 1727 1960
0 2147 6 1 2 1730 1961
0 2148 7 1 4 815 1267 363 67
0 2149 5 1 1 819
0 2150 7 1 2 822 831
0 2151 5 1 1 833
0 2152 5 1 1 823
0 2153 5 1 1 834
0 2154 7 1 2 824 837
0 2155 5 1 1 826
0 2156 5 1 1 838
0 2157 7 1 2 827 840
0 2158 9 16 1 847
0 2175 9 2 1 849
0 2178 6 1 2 1764 1981
0 2179 6 1 2 1766 1982
0 2180 5 1 1 841
0 2181 7 1 2 843 664
0 2183 5 1 1 844
0 2184 7 1 2 667 846
0 2185 6 2 2 677 859
0 2188 6 2 2 678 856
0 2191 6 2 2 673 860
0 2194 6 2 2 674 857
0 2197 6 2 2 680 853
0 2200 6 2 2 681 850
0 2203 6 2 2 675 855
0 2206 6 2 2 676 852
0 2209 5 1 1 862
0 2210 5 1 1 865
0 2211 7 1 2 863 866
0 2212 9 8 1 868
0 2221 9 8 1 869
0 2230 5 1 1 882
0 2231 5 1 1 884
0 2232 5 1 1 885
0 2233 5 1 1 887
0 2234 5 1 1 871
0 2235 5 1 1 872
0 2236 5 1 1 873
0 2237 5 1 1 875
0 2238 3 1 3 2022 1643 2023
0 2239 3 1 3 2024 1644 2025
0 2240 3 1 3 2026 1645 2027
0 2241 3 1 3 2028 1646 2029
0 2242 3 1 3 2030 1647 2031
0 2243 3 1 3 2032 1648 2033
0 2244 3 1 3 2034 1649 2035
0 2245 3 1 3 2036 1650 2037
0 2270 7 2 2 1986 1673
0 2277 7 2 2 1987 1675
0 2282 7 2 2 1988 1676
0 2287 7 2 2 1989 1677
0 2294 7 2 2 1990 1679
0 2299 7 2 2 1991 1680
0 2304 9 2 1 927
0 2307 7 2 2 942 351
0 2310 6 2 2 943 352
0 2313 9 2 1 811
0 2316 9 2 1 813
0 2319 9 2 1 812
0 2322 9 2 1 814
0 2325 6 2 2 1940 2133
0 2328 6 2 2 2134 2135
0 2331 6 2 2 2136 2137
0 2334 6 2 2 2138 2139
0 2341 6 1 2 949 2141
0 2342 6 1 2 946 2142
0 2347 7 1 2 412 2144
0 2348 7 1 3 2146 391 1726
0 2349 7 1 2 436 2147
0 2350 7 1 2 2148 633
0 2351 7 1 2 423 2150
0 2352 7 1 2 1735 2153
0 2353 7 1 2 447 2154
0 2354 7 1 2 1725 2156
0 2355 7 1 2 434 2157
0 2374 5 1 1 2178
0 2375 5 1 1 2179
0 2376 7 2 2 784 2180
0 2379 7 2 2 1721 2181
0 2398 7 1 2 364 2211
0 2417 7 1 3 974 231 1873
0 2418 7 1 3 975 275 648
0 2419 7 1 2 970 2238
0 2420 7 1 3 976 237 1878
0 2421 7 1 3 977 276 649
0 2422 7 1 2 971 2239
0 2425 7 1 3 978 243 1883
0 2426 7 1 3 979 277 650
0 2427 7 1 2 972 2240
0 2430 7 1 3 980 249 1888
0 2431 7 1 3 981 278 651
0 2432 7 1 2 973 2241
0 2435 7 1 3 960 256 1893
0 2436 7 1 3 961 279 660
0 2437 7 1 2 954 2242
0 2438 7 1 3 963 263 1898
0 2439 7 1 3 964 280 656
0 2440 7 1 2 955 2243
0 2443 7 1 3 966 269 1903
0 2444 7 1 3 967 281 657
0 2445 7 1 2 957 2244
0 2448 7 1 3 968 273 1908
0 2449 7 1 3 969 282 658
0 2450 7 1 2 958 2245
0 2467 5 1 1 1066
0 2468 5 1 1 1069
0 2469 5 1 1 1071
0 2470 5 1 1 1073
0 2471 6 2 2 2341 2342
0 2474 5 1 1 1075
0 2475 5 1 1 1077
0 2476 5 1 1 1079
0 2477 5 1 1 1081
0 2478 3 1 2 2348 1729
0 2481 5 1 1 1014
0 2482 7 1 2 1015 669
0 2483 7 2 2 2349 2183
0 2486 7 1 2 2374 1346
0 2487 7 1 2 2375 1350
0 2488 9 8 1 1016
0 2497 9 8 1 1018
0 2506 9 8 1 1020
0 2515 9 8 1 1022
0 2524 9 8 1 1024
0 2533 9 8 1 1026
0 2542 9 8 1 1028
0 2551 9 8 1 1030
0 2560 9 8 1 1017
0 2569 9 8 1 1019
0 2578 9 8 1 1021
0 2587 9 8 1 1023
0 2596 9 8 1 1025
0 2605 9 8 1 1027
0 2614 9 8 1 1029
0 2623 9 8 1 1031
0 2632 5 1 1 1032
0 2633 7 1 2 1033 888
0 2634 5 1 1 1034
0 2635 7 1 2 1035 893
0 2636 5 1 1 1036
0 2637 7 1 2 1037 894
0 2638 5 1 1 1038
0 2639 7 1 2 1039 897
0 2640 5 1 1 1040
0 2641 7 1 2 1041 876
0 2642 5 1 1 1042
0 2643 7 1 2 1043 878
0 2644 5 1 1 1044
0 2645 7 1 2 1045 879
0 2646 5 1 1 1046
0 2647 7 1 2 1047 881
0 2648 3 3 3 1048 898 982
0 2652 4 3 3 1049 899 983
0 2656 3 2 3 2417 2418 2419
0 2659 3 2 3 2420 2421 2422
0 2662 3 3 3 1050 902 986
0 2666 4 3 3 1051 903 987
0 2670 3 2 3 2425 2426 2427
0 2673 3 3 3 1052 904 988
0 2677 4 3 3 1053 905 989
0 2681 3 2 3 2430 2431 2432
0 2684 3 3 3 1054 906 990
0 2688 4 3 3 1055 907 991
0 2692 3 4 3 2435 2436 2437
0 2697 3 4 3 2438 2439 2440
0 2702 3 3 3 1056 910 994
0 2706 4 3 3 1057 911 995
0 2710 3 4 3 2443 2444 2445
0 2715 3 3 3 1058 912 996
0 2719 4 3 3 1059 918 997
0 2723 3 4 3 2448 2449 2450
0 2728 5 1 1 1060
0 2729 5 1 1 998
0 2730 7 1 2 797 999
0 2731 5 1 1 1000
0 2732 7 1 2 799 1001
0 2733 5 1 1 1002
0 2734 7 1 2 800 1003
0 2735 5 1 1 1004
0 2736 7 1 2 801 1005
0 2737 5 1 1 1006
0 2738 7 1 2 802 1007
0 2739 5 1 1 1008
0 2740 7 1 2 804 1009
0 2741 5 1 1 1010
0 2742 7 1 2 805 1011
0 2743 5 1 1 1012
0 2744 7 1 2 806 1013
0 2745 3 1 3 1083 951 1085
0 2746 4 1 3 1084 952 1086
0 2748 6 1 2 1070 2467
0 2749 6 1 2 1068 2468
0 2750 6 1 2 1074 2469
0 2751 6 1 2 1072 2470
0 2754 6 1 2 1078 2474
0 2755 6 1 2 1076 2475
0 2756 6 1 2 1082 2476
0 2757 6 1 2 1080 2477
0 2758 7 2 2 785 2481
0 2761 7 2 2 816 2482
0 2764 7 2 2 2478 1770
0 2768 3 1 3 2486 1789 1790
0 2769 3 1 3 2487 1797 1798
0 2898 7 1 2 365 2633
0 2899 7 1 2 376 2635
0 2900 7 1 2 381 2637
0 2901 7 1 2 394 2639
0 2962 5 1 1 2746
0 2966 6 1 2 2748 2749
0 2967 6 2 2 2750 2751
0 2970 9 2 1 1087
0 2973 6 3 2 2754 2755
0 2977 6 2 2 2756 2757
0 2980 7 1 2 1088 2143
0 2984 5 1 1 1091
0 2985 5 1 1 1099
0 2986 5 1 1 1107
0 2987 5 1 1 1115
0 2988 5 1 1 1124
0 2989 5 1 1 1132
0 2990 5 1 1 1140
0 2991 5 1 1 1148
0 2992 5 1 1 1092
0 2993 5 1 1 1100
0 2994 5 1 1 1108
0 2995 5 1 1 1116
0 2996 5 1 1 1125
0 2997 5 1 1 1133
0 2998 5 1 1 1141
0 2999 5 1 1 1149
0 3000 5 1 1 1093
0 3001 5 1 1 1101
0 3002 5 1 1 1109
0 3003 5 1 1 1118
0 3004 5 1 1 1126
0 3005 5 1 1 1134
0 3006 5 1 1 1142
0 3007 5 1 1 1150
0 3008 5 1 1 1094
0 3009 5 1 1 1102
0 3010 5 1 1 1110
0 3011 5 1 1 1119
0 3012 5 1 1 1127
0 3013 5 1 1 1135
0 3014 5 1 1 1143
0 3015 5 1 1 1151
0 3016 5 1 1 1095
0 3017 5 1 1 1103
0 3018 5 1 1 1111
0 3019 5 1 1 1120
0 3020 5 1 1 1128
0 3021 5 1 1 1136
0 3022 5 1 1 1144
0 3023 5 1 1 1152
0 3024 5 1 1 1096
0 3025 5 1 1 1104
0 3026 5 1 1 1112
0 3027 5 1 1 1121
0 3028 5 1 1 1129
0 3029 5 1 1 1137
0 3030 5 1 1 1145
0 3031 5 1 1 1153
0 3032 5 1 1 1097
0 3033 5 1 1 1105
0 3034 5 1 1 1113
0 3035 5 1 1 1122
0 3036 5 1 1 1130
0 3037 5 1 1 1138
0 3038 5 1 1 1146
0 3039 5 1 1 1154
0 3040 5 1 1 1098
0 3041 5 1 1 1106
0 3042 5 1 1 1114
0 3043 5 1 1 1123
0 3044 5 1 1 1131
0 3045 5 1 1 1139
0 3046 5 1 1 1147
0 3047 5 1 1 1155
0 3048 5 1 1 1156
0 3049 5 1 1 1164
0 3050 5 1 1 1172
0 3051 5 1 1 1181
0 3052 5 1 1 1189
0 3053 5 1 1 1199
0 3054 5 1 1 1208
0 3055 5 1 1 1216
0 3056 5 1 1 1157
0 3057 5 1 1 1165
0 3058 5 1 1 1173
0 3059 5 1 1 1182
0 3060 5 1 1 1190
0 3061 5 1 1 1200
0 3062 5 1 1 1209
0 3063 5 1 1 1217
0 3064 5 1 1 1158
0 3065 5 1 1 1166
0 3066 5 1 1 1174
0 3067 5 1 1 1183
0 3068 5 1 1 1191
0 3069 5 1 1 1201
0 3070 5 1 1 1210
0 3071 5 1 1 1218
0 3072 5 1 1 1159
0 3073 5 1 1 1167
0 3074 5 1 1 1175
0 3075 5 1 1 1184
0 3076 5 1 1 1192
0 3077 5 1 1 1203
0 3078 5 1 1 1211
0 3079 5 1 1 1220
0 3080 5 1 1 1160
0 3081 5 1 1 1168
0 3082 5 1 1 1176
0 3083 5 1 1 1185
0 3084 5 1 1 1193
0 3085 5 1 1 1204
0 3086 5 1 1 1212
0 3087 5 1 1 1221
0 3088 5 1 1 1161
0 3089 5 1 1 1169
0 3090 5 1 1 1177
0 3091 5 1 1 1186
0 3092 5 1 1 1194
0 3093 5 1 1 1205
0 3094 5 1 1 1213
0 3095 5 1 1 1222
0 3096 5 1 1 1162
0 3097 5 1 1 1170
0 3098 5 1 1 1178
0 3099 5 1 1 1187
0 3100 5 1 1 1195
0 3101 5 1 1 1206
0 3102 5 1 1 1214
0 3103 5 1 1 1223
0 3104 5 1 1 1163
0 3105 5 1 1 1171
0 3106 5 1 1 1180
0 3107 5 1 1 1188
0 3108 5 1 1 1198
0 3109 5 1 1 1207
0 3110 5 1 1 1215
0 3111 5 1 1 1224
0 3112 9 2 1 1231
0 3115 5 2 1 1232
0 3118 5 1 1 1228
0 3119 7 2 2 2768 1674
0 3122 9 2 1 1233
0 3125 5 2 1 1234
0 3128 9 2 1 1241
0 3131 5 2 1 1242
0 3134 5 1 1 1238
0 3135 9 2 1 1249
0 3138 5 2 1 1265
0 3141 5 1 1 1246
0 3142 9 2 1 1278
0 3145 5 2 1 1280
0 3148 5 1 1 1274
0 3149 7 2 2 2769 1678
0 3152 9 2 1 1283
0 3155 5 2 1 1284
0 3158 9 2 1 1293
0 3161 5 2 1 1294
0 3164 5 1 1 1290
0 3165 9 2 1 1305
0 3168 5 2 1 1307
0 3171 5 1 1 1301
0 3172 7 2 2 919 1225
0 3175 7 2 2 922 1235
0 3178 7 2 2 924 1243
0 3181 7 2 2 925 1266
0 3184 7 2 2 933 1287
0 3187 7 2 2 934 1297
0 3190 5 1 1 1281
0 3191 5 1 1 1285
0 3192 5 1 1 1295
0 3193 5 1 1 1308
0 3194 7 1 5 1282 1286 1296 1309 1459
3 3195 6 0 2 2745 2962
0 3196 5 1 1 2966
0 3206 3 1 3 2980 2145 2347
0 3207 7 1 2 124 2984
0 3208 7 1 2 161 2985
0 3209 7 1 2 152 2986
0 3210 7 1 2 144 2987
0 3211 7 1 2 138 2988
0 3212 7 1 2 133 2989
0 3213 7 1 2 129 2990
0 3214 7 1 2 126 2991
0 3215 7 1 2 127 2992
0 3216 7 1 2 355 2993
0 3217 7 1 2 162 2994
0 3218 7 1 2 153 2995
0 3219 7 1 2 145 2996
0 3220 7 1 2 139 2997
0 3221 7 1 2 134 2998
0 3222 7 1 2 130 2999
0 3223 7 1 2 131 3000
0 3224 7 1 2 367 3001
0 3225 7 1 2 356 3002
0 3226 7 1 2 163 3003
0 3227 7 1 2 154 3004
0 3228 7 1 2 146 3005
0 3229 7 1 2 140 3006
0 3230 7 1 2 135 3007
0 3231 7 1 2 136 3008
0 3232 7 1 2 383 3009
0 3233 7 1 2 368 3010
0 3234 7 1 2 357 3011
0 3235 7 1 2 164 3012
0 3236 7 1 2 155 3013
0 3237 7 1 2 147 3014
0 3238 7 1 2 141 3015
0 3239 7 1 2 142 3016
0 3240 7 1 2 396 3017
0 3241 7 1 2 384 3018
0 3242 7 1 2 369 3019
0 3243 7 1 2 358 3020
0 3244 7 1 2 165 3021
0 3245 7 1 2 156 3022
0 3246 7 1 2 148 3023
0 3247 7 1 2 149 3024
0 3248 7 1 2 404 3025
0 3249 7 1 2 397 3026
0 3250 7 1 2 385 3027
0 3251 7 1 2 370 3028
0 3252 7 1 2 359 3029
0 3253 7 1 2 166 3030
0 3254 7 1 2 157 3031
0 3255 7 1 2 158 3032
0 3256 7 1 2 414 3033
0 3257 7 1 2 405 3034
0 3258 7 1 2 398 3035
0 3259 7 1 2 386 3036
0 3260 7 1 2 371 3037
0 3261 7 1 2 360 3038
0 3262 7 1 2 167 3039
0 3263 7 1 2 168 3040
0 3264 7 1 2 425 3041
0 3265 7 1 2 415 3042
0 3266 7 1 2 406 3043
0 3267 7 1 2 399 3044
0 3268 7 1 2 387 3045
0 3269 7 1 2 372 3046
0 3270 7 1 2 361 3047
0 3271 7 1 2 286 3048
0 3272 7 1 2 373 3049
0 3273 7 1 2 388 3050
0 3274 7 1 2 400 3051
0 3275 7 1 2 407 3052
0 3276 7 1 2 416 3053
0 3277 7 1 2 426 3054
0 3278 7 1 2 437 3055
0 3279 7 1 2 296 3056
0 3280 7 1 2 389 3057
0 3281 7 1 2 401 3058
0 3282 7 1 2 408 3059
0 3283 7 1 2 417 3060
0 3284 7 1 2 427 3061
0 3285 7 1 2 438 3062
0 3286 7 1 2 287 3063
0 3287 7 1 2 305 3064
0 3288 7 1 2 402 3065
0 3289 7 1 2 409 3066
0 3290 7 1 2 418 3067
0 3291 7 1 2 428 3068
0 3292 7 1 2 439 3069
0 3293 7 1 2 288 3070
0 3294 7 1 2 297 3071
0 3295 7 1 2 312 3072
0 3296 7 1 2 410 3073
0 3297 7 1 2 419 3074
0 3298 7 1 2 429 3075
0 3299 7 1 2 440 3076
0 3300 7 1 2 289 3077
0 3301 7 1 2 298 3078
0 3302 7 1 2 306 3079
0 3303 7 1 2 318 3080
0 3304 7 1 2 420 3081
0 3305 7 1 2 430 3082
0 3306 7 1 2 441 3083
0 3307 7 1 2 290 3084
0 3308 7 1 2 299 3085
0 3309 7 1 2 307 3086
0 3310 7 1 2 313 3087
0 3311 7 1 2 323 3088
0 3312 7 1 2 431 3089
0 3313 7 1 2 442 3090
0 3314 7 1 2 291 3091
0 3315 7 1 2 300 3092
0 3316 7 1 2 308 3093
0 3317 7 1 2 314 3094
0 3318 7 1 2 319 3095
0 3319 7 1 2 327 3096
0 3320 7 1 2 443 3097
0 3321 7 1 2 292 3098
0 3322 7 1 2 301 3099
0 3323 7 1 2 309 3100
0 3324 7 1 2 315 3101
0 3325 7 1 2 320 3102
0 3326 7 1 2 324 3103
0 3327 7 1 2 329 3104
0 3328 7 1 2 293 3105
0 3329 7 1 2 302 3106
0 3330 7 1 2 310 3107
0 3331 7 1 2 316 3108
0 3332 7 1 2 321 3109
0 3333 7 1 2 325 3110
0 3334 7 1 2 328 3111
0 3383 7 1 5 3190 3191 3192 3193 555
0 3384 9 2 1 1326
0 3387 7 1 2 3196 1736
0 3388 7 1 2 1327 2149
0 3389 7 1 2 1321 1737
0 3390 4 1 8 3207 3208 3209 3210 3211 3212 3213 3214
0 3391 4 1 8 3215 3216 3217 3218 3219 3220 3221 3222
0 3392 4 1 8 3223 3224 3225 3226 3227 3228 3229 3230
0 3393 4 1 8 3231 3232 3233 3234 3235 3236 3237 3238
0 3394 4 1 8 3239 3240 3241 3242 3243 3244 3245 3246
0 3395 4 1 8 3247 3248 3249 3250 3251 3252 3253 3254
0 3396 4 1 8 3255 3256 3257 3258 3259 3260 3261 3262
0 3397 4 1 8 3263 3264 3265 3266 3267 3268 3269 3270
0 3398 4 1 8 3271 3272 3273 3274 3275 3276 3277 3278
0 3399 4 1 8 3279 3280 3281 3282 3283 3284 3285 3286
0 3400 4 1 8 3287 3288 3289 3290 3291 3292 3293 3294
0 3401 4 1 8 3295 3296 3297 3298 3299 3300 3301 3302
0 3402 4 1 8 3303 3304 3305 3306 3307 3308 3309 3310
0 3403 4 1 8 3311 3312 3313 3314 3315 3316 3317 3318
0 3404 4 1 8 3319 3320 3321 3322 3323 3324 3325 3326
0 3405 4 1 8 3327 3328 3329 3330 3331 3332 3333 3334
0 3406 7 1 2 3206 2641
0 3407 7 2 3 171 1226 1329
0 3410 7 2 3 182 1227 1332
0 3413 7 1 3 192 1229 1333
0 3414 7 1 3 205 1230 1330
0 3415 3 3 3 1335 900 984
0 3419 4 3 3 1336 901 985
0 3423 7 2 3 172 1236 1356
0 3426 7 2 3 183 1237 1359
0 3429 7 1 3 193 1239 1360
0 3430 7 1 3 206 1240 1357
0 3431 7 2 3 173 1244 1361
0 3434 7 2 3 184 1245 1364
0 3437 7 1 3 194 1247 1365
0 3438 7 1 3 207 1248 1362
0 3439 7 2 3 174 1269 1367
0 3442 7 2 3 185 1270 1370
0 3445 7 1 3 195 1275 1371
0 3446 7 1 3 208 1277 1368
0 3447 3 3 3 1372 908 992
0 3451 4 3 3 1373 909 993
0 3455 7 2 3 175 1288 1378
0 3458 7 2 3 186 1289 1380
0 3461 7 1 3 196 1291 1381
0 3462 7 1 3 209 1292 1379
0 3463 7 2 3 176 1299 1382
0 3466 7 2 3 187 1300 1385
0 3469 7 1 3 197 1303 1386
0 3470 7 1 3 210 1304 1383
0 3471 3 1 2 3194 3383
0 3472 9 2 1 1317
0 3475 9 2 1 1319
0 3478 9 2 1 1318
0 3481 9 2 1 1320
0 3484 9 2 1 1323
0 3487 9 2 1 1324
0 3490 9 2 1 1387
0 3493 9 2 1 1388
0 3496 9 2 1 1389
0 3499 9 2 1 1390
0 3502 9 2 1 1391
0 3505 9 2 1 1392
0 3508 9 2 1 1393
0 3511 9 2 1 1394
0 3514 9 2 1 1395
0 3517 9 2 1 1396
0 3520 9 2 1 1397
0 3523 9 2 1 1398
0 3534 4 1 2 3387 2350
0 3535 3 1 3 3388 2151 2351
0 3536 4 1 2 3389 1966
0 3537 7 1 2 3390 2209
0 3538 7 1 2 3398 2210
0 3539 7 1 2 3391 1842
0 3540 7 1 2 3399 696
0 3541 7 1 2 3392 1843
0 3542 7 1 2 3400 697
0 3543 7 1 2 3393 1844
0 3544 7 1 2 3401 698
0 3545 7 1 2 3394 1845
0 3546 7 1 2 3402 700
0 3547 7 1 2 3395 1846
0 3548 7 1 2 3403 701
0 3549 7 1 2 3396 1847
0 3550 7 1 2 3404 703
0 3551 7 1 2 3397 1848
0 3552 7 1 2 3405 704
0 3557 3 1 3 3413 3414 3118
0 3568 3 1 3 3429 3430 3134
0 3573 3 1 3 3437 3438 3141
0 3578 3 1 3 3445 3446 3148
0 3589 3 1 3 3461 3462 3164
0 3594 3 1 3 3469 3470 3171
0 3605 7 1 2 3471 2728
0 3626 5 1 1 1453
0 3627 5 1 1 1455
0 3628 5 1 1 1462
0 3629 5 1 1 1457
0 3630 5 1 1 1448
0 3631 5 1 1 1450
0 3632 7 1 2 3536 2152
0 3633 7 1 2 3534 2155
0 3634 3 1 3 3537 3538 2398
0 3635 3 1 2 3539 3540
0 3636 3 1 2 3541 3542
0 3637 3 1 2 3543 3544
0 3638 3 1 2 3545 3546
0 3639 3 1 2 3547 3548
0 3640 3 1 2 3549 3550
0 3641 3 1 2 3551 3552
0 3642 7 1 2 3535 2643
0 3643 3 1 2 1410 1412
0 3644 4 1 2 1411 1413
0 3645 7 2 3 177 1414 1341
0 3648 7 2 3 188 1415 1354
0 3651 7 1 3 198 1417 1355
0 3652 7 1 3 211 1418 1342
0 3653 5 1 1 1419
0 3654 3 2 2 1420 1422
0 3657 4 1 2 1421 1423
0 3658 3 2 2 1424 1428
0 3661 4 1 2 1425 1429
0 3662 3 1 2 1430 1432
0 3663 4 1 2 1431 1433
0 3664 7 2 3 178 1434 1374
0 3667 7 2 3 189 1435 1376
0 3670 7 1 3 199 1437 1377
0 3671 7 1 3 212 1438 1375
0 3672 5 1 1 1439
0 3673 3 2 2 1440 1442
0 3676 4 1 2 1441 1443
0 3677 3 2 2 1444 1446
0 3680 4 1 2 1445 1447
0 3681 5 1 1 1472
0 3682 7 2 2 921 1416
0 3685 5 1 1 1476
0 3686 5 1 1 1479
0 3687 5 1 1 1482
0 3688 5 1 1 1485
0 3689 5 1 1 1491
0 3690 7 2 2 936 1436
0 3693 5 1 1 1497
0 3694 5 1 1 1500
0 3695 5 1 1 1503
0 3696 5 1 1 1494
0 3697 9 2 1 1399
0 3700 9 2 1 1400
0 3703 5 1 1 1465
0 3704 5 1 1 1488
0 3705 6 1 2 1451 3630
0 3706 6 1 2 1449 3631
0 3707 6 1 2 1456 3626
0 3708 6 1 2 1454 3627
0 3711 3 1 3 3632 2352 2353
0 3712 3 1 3 3633 2354 2355
0 3713 7 1 2 3634 2632
0 3714 7 1 2 3635 2634
0 3715 7 1 2 3636 2636
0 3716 7 1 2 3637 2638
0 3717 7 1 2 3638 2640
0 3718 7 1 2 3639 2642
0 3719 7 1 2 3640 2644
0 3720 7 1 2 3641 2646
0 3721 7 5 2 3644 3557
0 3731 3 1 3 3651 3652 3653
0 3734 7 3 2 3657 3568
0 3740 7 2 2 3661 3573
0 3743 7 5 2 3663 3578
0 3753 3 1 3 3670 3671 3672
0 3756 7 3 2 3676 3589
0 3762 7 2 2 3680 3594
0 3765 5 1 1 3643
0 3766 5 1 1 3662
0 3773 6 1 2 3705 3706
0 3774 6 1 2 3707 3708
0 3775 6 1 2 1535 3628
0 3776 5 1 1 1536
0 3777 6 1 2 1533 3629
0 3778 5 1 1 1534
0 3779 7 1 2 3712 2645
0 3780 7 1 2 3711 2647
0 3786 3 2 2 1506 1514
0 3789 4 1 2 1513 1515
0 3800 3 2 2 1521 1523
0 3803 4 1 2 1522 1524
0 3809 7 2 2 1516 928
0 3812 7 2 2 1518 930
0 3815 7 2 2 1525 937
0 3818 7 2 2 1527 939
0 3821 9 2 1 1529
0 3824 9 2 1 1530
0 3827 9 2 1 1531
0 3830 9 2 1 1532
3 3833 6 0 2 3773 3774
0 3834 6 1 2 1463 3776
0 3835 6 1 2 1458 3778
0 3838 7 4 2 3789 3731
0 3845 7 4 2 3803 3753
0 3850 9 2 1 1537
0 3855 9 2 1 1542
0 3858 9 2 1 1545
0 3861 9 2 1 1547
0 3865 9 2 1 1552
0 3868 9 2 1 1555
0 3884 6 1 2 3775 3834
0 3885 6 1 2 3777 3835
0 3894 6 1 2 1538 1557
0 3895 6 1 2 1548 1559
0 3898 5 1 1 1570
0 3899 5 1 1 1572
0 3906 5 1 1 1576
0 3911 5 1 1 1574
0 3912 7 1 2 1558 1912
0 3913 9 2 1 1564
0 3916 7 1 2 1560 931
0 3917 9 2 1 1568
0 3920 5 1 1 1561
0 3921 9 2 1 1569
0 3924 5 1 1 3884
0 3925 5 1 1 3885
0 3926 7 3 4 1539 1578 1543 1546
0 3930 6 1 3 1540 1601 1517
0 3931 6 1 4 1519 1602 1544 1541
0 3932 7 2 4 1549 1604 1553 1556
0 3935 6 1 3 1550 1605 1526
0 3936 6 1 4 1528 1606 1554 1551
0 3937 9 2 1 1603
0 3940 9 2 1 1607
0 3947 5 1 1 3912
0 3948 5 1 1 3916
0 3950 9 2 1 1608
0 3953 9 2 1 1609
0 3956 9 2 1 1610
0 3959 9 2 1 1611
0 3962 9 2 1 1612
0 3965 9 2 1 1613
0 3968 9 2 1 1614
0 3971 9 2 1 1615
0 3974 9 2 1 1616
0 3977 9 2 1 1617
0 3980 9 2 1 1618
0 3983 9 2 1 1619
3 3987 6 0 2 3924 3925
0 3992 6 2 4 3765 3894 3930 3931
0 3996 6 2 4 3766 3895 3935 3936
0 4013 5 1 1 1624
3 4028 7 0 2 1629 1626
0 4029 6 1 2 1637 3681
0 4030 6 1 2 1641 3686
0 4031 6 1 2 1653 3688
0 4032 6 1 2 1657 3689
0 4033 6 1 2 1661 3693
0 4034 6 1 2 1665 3695
0 4035 9 2 1 1627
0 4042 5 1 1 1638
0 4043 5 1 1 1639
0 4044 6 1 2 1640 3685
0 4045 5 1 1 1642
0 4046 5 1 1 1651
0 4047 6 1 2 1652 3687
0 4048 5 1 1 1654
0 4049 5 1 1 1658
0 4050 5 1 1 1662
0 4051 5 1 1 1663
0 4052 6 1 2 1664 3694
0 4053 5 1 1 1666
0 4054 5 1 1 1659
0 4055 6 1 2 1660 3696
0 4056 7 1 2 1630 1061
0 4057 5 1 1 1635
0 4058 6 1 2 1636 3703
0 4059 9 2 1 1631
0 4062 9 2 1 1632
0 4065 5 1 1 1655
0 4066 6 1 2 1656 3704
0 4067 9 2 1 1633
0 4070 9 2 1 1634
0 4073 6 1 2 1628 1671
0 4074 5 1 1 1668
0 4075 6 1 2 1473 4042
0 4076 6 1 2 1480 4045
0 4077 6 1 2 1486 4048
0 4078 6 1 2 1492 4049
0 4079 6 1 2 1498 4050
0 4080 6 1 2 1504 4053
0 4085 6 1 2 1477 4043
0 4086 6 1 2 1483 4046
0 4088 6 1 2 1501 4051
0 4090 6 1 2 1495 4054
0 4091 7 2 2 1672 940
0 4094 3 3 2 3605 4056
0 4098 6 1 2 1466 4057
0 4101 6 1 2 1489 4065
0 4104 7 1 2 4073 4074
0 4105 6 1 2 4075 4029
0 4106 6 1 2 1685 3899
0 4107 6 1 2 4076 4030
0 4108 6 1 2 4077 4031
0 4109 6 1 2 4078 4032
0 4110 6 1 2 1689 3906
0 4111 6 1 2 4079 4033
0 4112 6 1 2 4080 4034
0 4113 5 1 1 1683
0 4114 6 1 2 1684 3898
0 4115 5 1 1 1686
0 4116 6 2 2 4085 4044
0 4119 6 2 2 4086 4047
0 4122 5 1 1 1690
0 4123 6 2 2 4088 4052
0 4126 5 1 1 1687
0 4127 6 1 2 1688 3911
0 4128 6 5 2 4090 4055
0 4139 6 2 2 4098 4058
0 4142 6 2 2 4101 4066
3 4145 5 0 1 4104
0 4146 5 1 1 4105
0 4147 6 1 2 1573 4115
0 4148 5 1 1 4107
0 4149 5 1 1 4108
0 4150 5 1 1 4109
0 4151 6 1 2 1577 4122
0 4152 5 1 1 4111
0 4153 5 1 1 4112
0 4154 6 1 2 1571 4113
0 4161 6 1 2 1575 4126
0 4167 9 6 1 1695
0 4174 9 4 1 1697
0 4182 9 2 1 1696
0 4186 7 2 2 332 1698
0 4189 7 1 2 4146 2230
0 4190 6 1 2 4147 4106
0 4191 7 1 2 4148 2232
0 4192 7 1 2 4149 2233
0 4193 7 1 2 4150 2234
0 4194 6 1 2 4151 4110
0 4195 7 1 2 4152 2236
0 4196 7 1 2 4153 2237
0 4197 6 2 2 4154 4114
0 4200 9 2 1 1700
0 4203 9 5 1 1701
0 4209 9 3 1 1702
0 4213 9 4 1 1703
0 4218 6 4 2 4161 4127
0 4223 9 4 1 1704
0 4238 7 1 2 1706 1622
0 4239 5 1 1 1711
0 4241 5 1 1 1716
0 4242 7 2 2 333 1705
0 4247 9 2 1 1707
0 4251 4 1 3 3713 4189 2898
0 4252 5 1 1 4190
0 4253 4 1 3 3715 4191 2900
0 4254 4 1 3 3716 4192 2901
0 4255 4 1 3 3717 4193 3406
0 4256 5 1 1 4194
0 4257 4 1 3 3719 4195 3779
0 4258 4 1 3 3720 4196 3780
0 4283 7 1 2 1719 1681
0 4284 7 2 2 1734 1682
0 4287 3 3 2 1566 4238
0 4291 5 1 1 1744
0 4295 5 1 1 1720
0 4296 9 2 1 1723
0 4299 5 1 1 1742
0 4303 7 1 2 4252 2231
0 4304 7 1 2 4256 2235
0 4305 9 4 1 1746
0 4310 3 3 2 1669 4283
0 4316 7 1 3 1739 1760 1751
0 4317 7 1 2 1740 1757
0 4318 7 1 3 1776 1708 1772
0 4319 7 2 2 1777 1709
0 4322 7 1 2 1724 1758
0 4325 6 1 2 1752 1620
0 4326 6 1 3 1753 1762 1732
0 4327 6 1 2 1773 1567
0 4328 6 1 3 1774 1710 1623
0 4329 6 1 2 1782 4013
0 4330 5 1 1 1783
0 4331 7 2 3 334 1699 4295
0 4335 7 2 2 4251 2730
0 4338 7 2 2 4253 2734
0 4341 7 2 2 4254 2736
0 4344 7 2 2 4255 2738
0 4347 7 2 2 4257 2742
0 4350 7 2 2 4258 2744
0 4353 9 2 1 1748
0 4356 9 2 1 1754
0 4359 9 2 1 1759
0 4362 9 2 1 1775
0 4365 9 2 1 1780
0 4368 9 2 1 1781
0 4371 7 2 2 1778 1778
0 4376 4 1 3 3714 4303 2899
0 4377 4 1 3 3718 4304 3642
0 4387 7 2 2 335 4317
0 4390 7 2 2 336 4318
0 4393 6 1 2 1625 4330
0 4398 9 2 1 1786
0 4413 9 2 1 1784
0 4416 6 2 3 3920 4325 4326
0 4421 3 2 2 1565 4322
0 4427 6 2 3 3948 4327 4328
0 4430 9 2 1 1804
0 4435 7 2 2 337 4316
0 4442 3 1 2 1823 1807
0 4443 7 2 4 1741 1810 1755 1763
0 4446 6 1 2 1811 1563
0 4447 6 1 3 1813 1749 1621
0 4448 6 1 4 1814 1750 1771 1733
0 4452 5 1 1 1841
0 4458 6 2 2 4329 4393
0 4461 5 1 1 1872
0 4462 5 1 1 1877
0 4463 6 1 2 1882 1460
0 4464 5 1 1 1886
0 4465 9 2 1 1816
0 4468 4 2 2 1825 1808
0 4472 7 2 2 4376 2732
0 4475 7 2 2 4377 2740
0 4479 9 2 1 1817
0 4484 5 1 1 1839
0 4486 5 1 1 1866
0 4487 6 1 2 1867 4299
0 4491 5 1 1 1868
0 4493 7 2 2 338 1820
0 4496 5 1 1 1897
0 4497 7 1 2 1805 1901
0 4498 7 2 2 4442 1769
0 4503 6 2 4 3947 4446 4447 4448
0 4506 5 1 1 1902
0 4507 5 1 1 1920
0 4508 5 1 1 1911
0 4509 6 1 2 1914 4452
0 4510 5 1 1 1915
0 4511 6 1 2 1916 4241
0 4515 6 1 2 587 4464
0 4526 5 1 1 1907
0 4527 6 1 2 1910 4484
0 4528 6 1 2 1743 4486
0 4529 5 1 1 1918
0 4530 6 1 2 1919 4491
0 4531 9 2 1 1887
0 4534 9 2 1 1891
0 4537 9 2 1 1892
0 4540 9 2 1 1896
0 4545 7 1 3 339 1822 4496
0 4549 7 2 2 340 1923
0 4552 6 1 2 1865 4508
0 4555 6 1 2 1717 4510
0 4558 5 1 1 1950
0 4559 6 2 2 4463 4515
0 4562 5 1 1 1928
0 4563 7 1 2 1819 1929
0 4564 9 3 1 1931
0 4568 5 1 1 1948
0 4569 9 2 1 1924
0 4572 6 1 2 1840 4526
0 4573 6 1 2 1871 4529
0 4576 6 2 2 4487 4528
0 4581 9 2 1 1925
0 4584 9 2 1 1927
0 4587 3 1 3 1310 1952 1312
0 4588 4 1 3 1311 1953 1313
3 4589 3 0 2 4545 4497
0 4593 6 2 2 4552 4509
0 4596 5 1 1 1956
0 4597 5 1 1 1958
0 4599 6 2 2 4555 4511
0 4602 5 1 1 1962
0 4603 5 1 1 1964
0 4608 7 1 3 341 1785 4562
0 4613 9 2 1 1954
0 4616 9 2 1 1955
0 4619 6 2 2 4572 4527
0 4623 6 2 2 4573 4530
0 4628 5 1 1 4588
0 4629 6 1 2 1974 4506
0 4630 5 1 1 1975
0 4635 5 1 1 1976
0 4636 6 1 2 1977 4291
0 4640 5 1 1 1978
0 4641 6 1 2 1979 4461
0 4642 5 1 1 1980
0 4643 6 1 2 1984 4462
0 4644 4 2 2 4608 4563
0 4647 7 2 2 1969 2128
0 4650 7 2 2 1970 2743
0 4656 9 2 1 1967
0 4659 9 2 1 1968
0 4664 9 2 1 1971
3 4667 7 0 2 4587 4628
0 4668 6 1 2 1906 4630
0 4669 5 1 1 1997
0 4670 6 1 2 1998 4239
0 4673 5 1 1 1999
0 4674 6 1 2 2000 4507
0 4675 6 1 2 1745 4635
0 4676 5 1 1 2001
0 4677 6 1 2 2002 4558
0 4678 6 1 2 1876 4640
0 4679 6 1 2 1881 4642
0 4687 5 1 1 1995
0 4688 6 1 2 1996 4568
0 4691 9 2 1 1985
0 4694 9 2 1 1992
0 4697 9 2 1 1993
0 4700 9 2 1 1994
0 4704 6 1 2 4629 4668
0 4705 6 1 2 1712 4669
0 4706 5 1 1 2009
0 4707 5 1 1 2011
0 4708 6 1 2 1921 4673
0 4711 6 2 2 4675 4636
0 4716 6 1 2 1951 4676
0 4717 6 3 2 4678 4641
0 4721 6 1 2 4679 4643
0 4722 9 3 1 2003
0 4726 5 1 1 2013
0 4727 3 2 3 2005 2007 1837
0 4730 4 2 3 2006 2008 1838
0 4733 6 1 2 1949 4687
0 4740 6 2 2 4705 4670
0 4743 6 3 2 4708 4674
0 4747 5 1 1 2015
0 4748 6 1 2 2016 4596
0 4749 5 1 1 2017
0 4750 6 1 2 2018 4597
0 4753 5 1 1 2019
0 4754 6 1 2 2020 4602
0 4755 5 1 1 2021
0 4756 6 1 2 2039 4603
0 4757 6 3 2 4716 4677
0 4769 6 2 2 4733 4688
0 4772 7 2 2 342 4704
0 4775 5 2 1 4721
0 4778 5 1 1 2051
0 4786 6 1 2 1957 4747
0 4787 6 1 2 1959 4749
0 4788 6 1 2 1963 4753
0 4789 6 1 2 1965 4755
0 4794 7 2 2 2040 2124
0 4797 7 2 2 2041 2735
0 4800 7 2 2 2042 2127
0 4805 9 2 1 2046
0 4808 7 2 2 2044 1932
0 4812 9 2 1 2049
3 4815 7 0 2 2050 4778
0 4816 5 1 1 2063
0 4817 5 1 1 2065
0 4818 6 3 2 4786 4748
0 4822 6 1 2 4787 4750
0 4823 6 2 2 4788 4754
0 4826 6 1 2 4789 4756
0 4829 6 1 2 2067 4726
0 4830 5 1 1 2069
0 4831 7 2 2 2056 2122
0 4838 7 2 2 2060 2126
0 4844 9 2 1 2054
0 4847 9 2 1 2055
0 4850 9 2 1 2058
0 4854 9 2 1 2061
0 4859 6 1 2 2066 4816
0 4860 6 1 2 2064 4817
0 4868 5 1 1 4826
0 4870 5 1 1 2077
0 4872 5 1 1 2080
0 4873 6 1 2 2014 4830
0 4876 3 3 3 2070 2072 1830
0 4880 4 2 3 2071 2074 1831
0 4885 5 1 1 2082
0 4889 5 2 1 4822
0 4895 6 1 2 4859 4860
0 4896 5 1 1 2096
0 4897 6 1 2 2097 4706
0 4898 5 1 1 2099
0 4899 6 1 2 2100 4707
0 4900 4 1 2 4868 1972
0 4901 7 1 4 2045 2062 2089 1973
0 4902 5 1 1 2101
0 4904 5 1 1 2104
0 4905 6 1 2 2105 4872
0 4906 6 1 2 4873 4829
0 4907 7 2 2 2085 2123
0 4913 7 2 2 2090 2125
0 4916 7 2 2 2086 2004
0 4920 5 1 1 2109
0 4921 7 2 2 4895 2184
0 4924 6 1 2 2010 4896
0 4925 6 1 2 2012 4898
0 4926 3 1 2 4900 4901
0 4928 6 1 2 2111 4870
0 4929 5 1 1 2112
0 4930 6 1 2 2081 4904
0 4931 5 1 1 4906
0 4937 9 2 1 2106
0 4940 9 2 1 2107
3 4944 7 0 2 2108 4920
0 4946 6 2 2 4924 4897
0 4949 6 1 2 4925 4899
0 4950 6 1 2 2117 4902
0 4951 5 1 1 2118
0 4952 6 1 2 2079 4929
0 4953 6 1 2 4930 4905
0 4954 7 2 2 4926 2737
0 4957 7 2 2 4931 2741
0 4964 3 1 3 1314 1089 2119
0 4965 4 1 3 1316 1090 2120
0 4968 5 1 1 4949
0 4969 6 1 2 2102 4951
0 4970 6 1 2 4952 4928
0 4973 7 2 2 4953 2739
0 4978 5 1 1 2129
0 4979 5 1 1 2131
0 4980 5 1 1 4965
0 4981 4 1 2 4968 2047
0 4982 7 1 4 2087 2059 2140 2048
0 4983 6 1 2 4950 4969
0 4984 5 1 1 4970
0 4985 7 2 2 2159 2121
0 4988 3 2 3 2115 2160 1832
0 4991 4 2 3 2116 2161 1834
0 4996 3 2 3 2075 2162 1835
0 4999 4 2 3 2076 2163 1836
3 5002 7 0 2 4964 4980
0 5007 3 1 2 4981 4982
0 5010 7 2 2 4983 2731
0 5013 7 2 2 4984 2733
0 5018 3 2 3 2094 2164 1937
0 5021 4 2 3 2095 2165 1938
0 5026 5 1 1 2170
0 5029 5 1 1 2174
0 5030 7 2 2 5007 2729
0 5039 9 2 1 2172
0 5042 9 2 1 2168
3 5045 7 0 2 2169 5026
0 5046 5 1 1 2192
3 5047 7 0 2 2173 5029
0 5050 3 4 3 2091 2177 1934
0 5055 4 2 3 2092 2182 1935
0 5058 3 2 3 2113 2186 1828
0 5061 4 2 3 2114 2187 1829
0 5066 7 2 4 2053 2176 2193 2171
0 5070 9 2 1 2189
3 5078 7 0 2 2190 5046
0 5080 3 4 3 2166 2195 1826
0 5085 4 2 3 2167 2196 1827
0 5094 6 1 2 2198 4885
0 5095 5 1 1 2199
0 5097 5 1 1 2201
3 5102 7 0 2 2204 2204
0 5103 5 1 1 2217
0 5108 6 1 2 2084 5095
0 5109 5 1 1 2222
0 5110 6 1 2 2223 5097
0 5111 9 2 1 2215
0 5114 7 2 2 2207 750
0 5117 9 2 1 2208
3 5120 7 0 2 2224 2224
3 5121 7 0 2 2216 5103
0 5122 6 2 2 5094 5108
0 5125 6 1 2 2202 5109
0 5128 7 2 2 751 2226
0 5133 7 2 4 2110 2218 2213 2228
0 5136 7 1 3 2214 2229 754
0 5139 9 2 1 2227
0 5145 6 2 2 5125 5110
0 5151 9 2 1 2246
0 5154 9 2 1 2247
0 5159 5 1 1 2250
0 5160 9 2 1 2248
0 5163 9 2 1 2249
0 5166 7 1 2 2219 2256
0 5173 7 1 2 2220 2257
0 5174 9 2 1 2252
0 5177 9 2 1 2253
0 5182 5 1 1 2258
0 5183 6 1 2 2259 5159
0 5184 9 2 1 2254
0 5188 9 2 1 2255
3 5192 5 0 1 5166
0 5193 4 1 2 5136 5173
0 5196 6 1 2 2262 4978
0 5197 5 1 1 2263
0 5198 6 1 2 2264 4979
0 5199 5 1 1 2265
0 5201 5 1 1 2266
0 5203 5 1 1 2268
0 5205 9 2 1 2260
0 5209 9 2 1 2261
0 5212 6 1 2 2251 5182
0 5215 7 1 2 221 5193
0 5217 5 1 1 2271
0 5219 5 1 1 2273
0 5220 6 1 2 2130 5197
0 5221 6 1 2 2132 5199
0 5222 5 1 1 2275
0 5223 6 1 2 2276 5201
0 5224 6 1 2 2278 5203
0 5225 5 1 1 2279
0 5228 6 2 2 5183 5212
3 5231 5 0 1 5215
0 5232 6 1 2 2280 5217
0 5233 5 1 1 2281
0 5234 6 1 2 2283 5219
0 5235 5 1 1 2284
0 5236 6 3 2 5196 5220
0 5240 6 1 2 5198 5221
0 5242 6 1 2 2267 5222
0 5243 6 1 2 2269 5225
0 5245 6 1 2 2272 5233
0 5246 6 1 2 2274 5235
0 5250 5 2 1 5240
0 5253 5 1 1 2285
0 5254 6 2 2 5242 5223
0 5257 6 1 2 5243 5224
0 5258 6 2 2 5232 5245
0 5261 6 1 2 5234 5246
0 5266 5 2 1 5257
0 5269 9 2 1 2288
0 5277 7 1 3 2289 2293 1062
0 5278 7 1 3 2291 2295 1064
0 5279 5 2 1 5261
0 5283 5 1 1 2301
0 5284 6 1 2 2302 5253
0 5285 7 1 3 2290 2298 1065
0 5286 7 1 3 2292 2300 1063
0 5289 9 2 1 2296
0 5292 9 2 1 2297
0 5295 6 1 2 2286 5283
0 5298 3 2 4 5277 5285 5278 5286
0 5303 9 2 1 2303
0 5306 9 2 1 2305
0 5309 6 2 2 5295 5284
0 5312 5 1 1 2309
0 5313 5 1 1 2306
0 5322 5 1 1 2318
0 5323 5 1 1 2315
0 5324 9 2 1 2312
0 5327 9 2 1 2314
0 5332 9 2 1 2321
0 5335 9 2 1 2323
0 5340 6 1 2 2324 5323
0 5341 6 1 2 2327 5322
0 5344 5 1 1 2329
0 5345 5 1 1 2326
0 5348 6 1 2 2330 5313
0 5349 6 1 2 2333 5312
0 5350 6 1 2 2317 5345
0 5351 6 1 2 2320 5344
0 5352 5 1 1 2335
0 5353 5 1 1 2332
0 5354 6 1 2 2308 5353
0 5355 6 1 2 2311 5352
0 5356 6 1 2 5350 5340
0 5357 6 1 2 5351 5341
0 5358 6 1 2 5348 5354
0 5359 6 1 2 5349 5355
3 5360 7 0 2 5356 5357
3 5361 6 0 2 5358 5359
2 2 1 1
2 3 1 1
2 4 1 1
2 5 1 1
2 6 1 1
2 7 1 1
2 8 1 1
2 9 1 1
2 10 1 1
2 11 1 1
2 12 1 1
2 14 1 13
2 15 1 13
2 16 1 13
2 17 1 13
2 18 1 13
2 19 1 13
2 21 1 20
2 22 1 20
2 23 1 20
2 24 1 20
2 25 1 20
2 26 1 20
2 27 1 20
2 28 1 20
2 29 1 20
2 30 1 20
2 31 1 20
2 32 1 20
2 34 1 33
2 35 1 33
2 36 1 33
2 37 1 33
2 38 1 33
2 39 1 33
2 40 1 33
2 42 1 41
2 43 1 41
2 44 1 41
2 46 1 45
2 47 1 45
2 48 1 45
2 49 1 45
2 51 1 50
2 52 1 50
2 53 1 50
2 54 1 50
2 55 1 50
2 56 1 50
2 57 1 50
2 59 1 58
2 60 1 58
2 61 1 58
2 62 1 58
2 63 1 58
2 64 1 58
2 65 1 58
2 66 1 58
2 67 1 58
2 69 1 68
2 70 1 68
2 71 1 68
2 72 1 68
2 73 1 68
2 74 1 68
2 75 1 68
2 76 1 68
2 78 1 77
2 79 1 77
2 80 1 77
2 81 1 77
2 82 1 77
2 83 1 77
2 84 1 77
2 85 1 77
2 86 1 77
2 88 1 87
2 89 1 87
2 90 1 87
2 91 1 87
2 92 1 87
2 93 1 87
2 94 1 87
2 95 1 87
2 96 1 87
2 98 1 97
2 99 1 97
2 100 1 97
2 101 1 97
2 102 1 97
2 103 1 97
2 104 1 97
2 105 1 97
2 106 1 97
2 108 1 107
2 109 1 107
2 110 1 107
2 111 1 107
2 112 1 107
2 113 1 107
2 114 1 107
2 115 1 107
2 117 1 116
2 118 1 116
2 119 1 116
2 120 1 116
2 121 1 116
2 122 1 116
2 123 1 116
2 126 1 125
2 127 1 125
2 129 1 128
2 130 1 128
2 131 1 128
2 133 1 132
2 134 1 132
2 135 1 132
2 136 1 132
2 138 1 137
2 139 1 137
2 140 1 137
2 141 1 137
2 142 1 137
2 144 1 143
2 145 1 143
2 146 1 143
2 147 1 143
2 148 1 143
2 149 1 143
2 151 1 150
2 152 1 150
2 153 1 150
2 154 1 150
2 155 1 150
2 156 1 150
2 157 1 150
2 158 1 150
2 160 1 159
2 161 1 159
2 162 1 159
2 163 1 159
2 164 1 159
2 165 1 159
2 166 1 159
2 167 1 159
2 168 1 159
2 170 1 169
2 171 1 169
2 172 1 169
2 173 1 169
2 174 1 169
2 175 1 169
2 176 1 169
2 177 1 169
2 178 1 169
2 180 1 179
2 181 1 179
2 182 1 179
2 183 1 179
2 184 1 179
2 185 1 179
2 186 1 179
2 187 1 179
2 188 1 179
2 189 1 179
2 191 1 190
2 192 1 190
2 193 1 190
2 194 1 190
2 195 1 190
2 196 1 190
2 197 1 190
2 198 1 190
2 199 1 190
2 201 1 200
2 202 1 200
2 203 1 200
2 204 1 200
2 205 1 200
2 206 1 200
2 207 1 200
2 208 1 200
2 209 1 200
2 210 1 200
2 211 1 200
2 212 1 200
2 214 1 213
2 215 1 213
2 216 1 213
2 217 1 213
2 218 1 213
2 219 1 213
2 220 1 213
2 221 1 213
2 224 1 223
2 225 1 223
2 227 1 226
2 228 1 226
2 229 1 226
2 230 1 226
2 231 1 226
2 233 1 232
2 234 1 232
2 235 1 232
2 236 1 232
2 237 1 232
2 239 1 238
2 240 1 238
2 241 1 238
2 242 1 238
2 243 1 238
2 245 1 244
2 246 1 244
2 247 1 244
2 248 1 244
2 249 1 244
2 251 1 250
2 252 1 250
2 253 1 250
2 254 1 250
2 255 1 250
2 256 1 250
2 258 1 257
2 259 1 257
2 260 1 257
2 261 1 257
2 262 1 257
2 263 1 257
2 265 1 264
2 266 1 264
2 267 1 264
2 268 1 264
2 269 1 264
2 271 1 270
2 272 1 270
2 273 1 270
2 275 1 274
2 276 1 274
2 277 1 274
2 278 1 274
2 279 1 274
2 280 1 274
2 281 1 274
2 282 1 274
2 284 1 283
2 285 1 283
2 286 1 283
2 287 1 283
2 288 1 283
2 289 1 283
2 290 1 283
2 291 1 283
2 292 1 283
2 293 1 283
2 295 1 294
2 296 1 294
2 297 1 294
2 298 1 294
2 299 1 294
2 300 1 294
2 301 1 294
2 302 1 294
2 304 1 303
2 305 1 303
2 306 1 303
2 307 1 303
2 308 1 303
2 309 1 303
2 310 1 303
2 312 1 311
2 313 1 311
2 314 1 311
2 315 1 311
2 316 1 311
2 318 1 317
2 319 1 317
2 320 1 317
2 321 1 317
2 323 1 322
2 324 1 322
2 325 1 322
2 327 1 326
2 328 1 326
2 331 1 330
2 332 1 330
2 333 1 330
2 334 1 330
2 335 1 330
2 336 1 330
2 337 1 330
2 338 1 330
2 339 1 330
2 340 1 330
2 341 1 330
2 342 1 330
2 344 1 343
2 345 1 343
2 346 1 343
2 347 1 343
2 348 1 343
2 351 1 350
2 352 1 350
2 353 1 655
2 354 1 655
2 355 1 655
2 356 1 655
2 357 1 655
2 358 1 655
2 359 1 655
2 360 1 655
2 361 1 655
2 362 1 665
2 363 1 665
2 364 1 665
2 365 1 665
2 366 1 670
2 367 1 670
2 368 1 670
2 369 1 670
2 370 1 670
2 371 1 670
2 372 1 670
2 373 1 670
2 374 1 679
2 375 1 679
2 376 1 679
2 377 1 683
2 378 1 683
2 379 1 686
2 380 1 686
2 381 1 686
2 382 1 690
2 383 1 690
2 384 1 690
2 385 1 690
2 386 1 690
2 387 1 690
2 388 1 690
2 389 1 690
2 390 1 699
2 391 1 699
2 392 1 702
2 393 1 702
2 394 1 702
2 395 1 706
2 396 1 706
2 397 1 706
2 398 1 706
2 399 1 706
2 400 1 706
2 401 1 706
2 402 1 706
2 403 1 715
2 404 1 715
2 405 1 715
2 406 1 715
2 407 1 715
2 408 1 715
2 409 1 715
2 410 1 715
2 411 1 724
2 412 1 724
2 413 1 727
2 414 1 727
2 415 1 727
2 416 1 727
2 417 1 727
2 418 1 727
2 419 1 727
2 420 1 727
2 421 1 736
2 422 1 736
2 423 1 736
2 424 1 740
2 425 1 740
2 426 1 740
2 427 1 740
2 428 1 740
2 429 1 740
2 430 1 740
2 431 1 740
2 432 1 749
2 433 1 749
2 434 1 749
2 435 1 753
2 436 1 753
2 437 1 753
2 438 1 753
2 439 1 753
2 440 1 753
2 441 1 753
2 442 1 753
2 443 1 753
2 444 1 763
2 445 1 763
2 446 1 763
2 447 1 763
2 448 1 769
2 449 1 769
2 450 1 772
2 451 1 772
2 452 1 772
2 453 1 772
2 454 1 772
2 455 1 772
2 456 1 779
2 457 1 779
2 458 1 782
2 459 1 782
2 460 1 782
2 461 1 786
2 462 1 786
2 463 1 786
2 464 1 786
2 465 1 786
2 466 1 786
2 467 1 794
2 468 1 794
2 469 1 794
2 470 1 798
2 471 1 798
2 472 1 798
2 473 1 798
2 474 1 803
2 475 1 803
2 476 1 803
2 477 1 803
2 478 1 803
2 479 1 803
2 480 1 803
2 481 1 803
2 482 1 803
2 483 1 803
2 484 1 803
2 485 1 803
2 486 1 803
2 487 1 803
2 488 1 803
2 489 1 803
2 490 1 821
2 491 1 821
2 492 1 821
2 493 1 825
2 494 1 825
2 495 1 825
2 496 1 829
2 497 1 829
2 498 1 832
2 499 1 832
2 500 1 836
2 501 1 836
2 502 1 839
2 503 1 839
2 504 1 842
2 505 1 842
2 506 1 845
2 507 1 845
2 508 1 848
2 509 1 848
2 510 1 851
2 511 1 851
2 512 1 854
2 513 1 854
2 514 1 854
2 515 1 858
2 516 1 858
2 517 1 861
2 518 1 861
2 519 1 864
2 520 1 864
2 521 1 867
2 522 1 867
2 523 1 870
2 524 1 870
2 525 1 870
2 526 1 874
2 527 1 874
2 528 1 877
2 529 1 877
2 530 1 880
2 531 1 880
2 532 1 883
2 533 1 883
2 534 1 886
2 535 1 886
2 536 1 892
2 537 1 892
2 538 1 896
2 539 1 896
2 540 1 896
2 541 1 896
2 542 1 896
2 543 1 896
2 544 1 896
2 545 1 896
2 546 1 896
2 547 1 896
2 548 1 896
2 549 1 896
2 550 1 896
2 551 1 896
2 552 1 896
2 553 1 896
2 554 1 917
2 555 1 917
2 556 1 920
2 557 1 920
2 558 1 923
2 559 1 923
2 560 1 926
2 561 1 926
2 562 1 929
2 563 1 929
2 564 1 932
2 565 1 932
2 566 1 935
2 567 1 935
2 568 1 938
2 569 1 938
2 570 1 941
2 571 1 941
2 572 1 944
2 573 1 944
2 574 1 947
2 575 1 947
2 576 1 950
2 577 1 950
2 578 1 953
2 579 1 953
2 580 1 956
2 581 1 956
2 582 1 959
2 583 1 959
2 584 1 962
2 585 1 962
2 586 1 965
2 587 1 965
2 588 1 1117
2 589 1 1117
2 590 1 1117
2 591 1 1117
2 592 1 1117
2 593 1 1117
2 594 1 1117
2 595 1 1117
2 596 1 1117
2 597 1 1117
2 598 1 1117
2 599 1 1117
2 600 1 1117
2 601 1 1117
2 602 1 1117
2 603 1 1117
2 604 1 1197
2 605 1 1197
2 606 1 1197
2 607 1 1197
2 608 1 1202
2 609 1 1202
2 610 1 1202
2 611 1 1202
2 612 1 1202
2 613 1 1202
2 614 1 1202
2 615 1 1202
2 616 1 1202
2 617 1 1202
2 618 1 1202
2 619 1 1202
2 620 1 1202
2 621 1 1202
2 622 1 1202
2 623 1 1202
2 624 1 1219
2 625 1 1219
2 626 1 1219
2 627 1 1219
2 628 1 1264
2 629 1 1264
2 630 1 1268
2 631 1 1268
2 632 1 1273
2 633 1 1273
2 634 1 1276
2 635 1 1276
2 636 1 1279
2 637 1 1279
2 638 1 1298
2 639 1 1298
2 640 1 1298
2 641 1 1302
2 642 1 1302
2 643 1 1302
2 644 1 1306
2 645 1 1306
2 646 1 1306
2 647 1 1306
2 648 1 1306
2 649 1 1306
2 650 1 1306
2 651 1 1306
2 652 1 1315
2 653 1 1315
2 654 1 1315
2 656 1 1315
2 657 1 1315
2 658 1 1315
2 659 1 1322
2 660 1 1322
2 661 1 1325
2 662 1 1325
2 663 1 1328
2 664 1 1328
2 666 1 1331
2 667 1 1331
2 668 1 1334
2 669 1 1334
2 671 1 1340
2 672 1 1340
2 673 1 1353
2 674 1 1353
2 675 1 1353
2 676 1 1353
2 677 1 1358
2 678 1 1358
2 680 1 1358
2 681 1 1358
2 682 1 1363
2 684 1 1363
2 685 1 1366
2 687 1 1366
2 688 1 1369
2 689 1 1369
2 691 1 1369
2 692 1 1369
2 693 1 1369
2 694 1 1369
2 695 1 1369
2 696 1 1369
2 697 1 1369
2 698 1 1369
2 700 1 1369
2 701 1 1369
2 703 1 1369
2 704 1 1369
2 705 1 1384
2 707 1 1384
2 708 1 1384
2 709 1 1384
2 710 1 1384
2 711 1 1384
2 712 1 1384
2 713 1 1384
2 714 1 1384
2 716 1 1384
2 717 1 1384
2 718 1 1384
2 719 1 1384
2 720 1 1384
2 721 1 1384
2 722 1 1384
2 723 1 1409
2 725 1 1409
2 726 1 1409
2 728 1 1409
2 729 1 1409
2 730 1 1409
2 731 1 1409
2 732 1 1409
2 733 1 1409
2 734 1 1409
2 735 1 1409
2 737 1 1409
2 738 1 1409
2 739 1 1409
2 741 1 1409
2 742 1 1409
2 743 1 1452
2 744 1 1452
2 745 1 1452
2 746 1 1452
2 747 1 1452
2 748 1 1452
2 750 1 1461
2 751 1 1461
2 752 1 1464
2 754 1 1464
2 755 1 1471
2 756 1 1471
2 757 1 1475
2 758 1 1475
2 759 1 1478
2 760 1 1478
2 761 1 1481
2 762 1 1481
2 764 1 1484
2 765 1 1484
2 766 1 1487
2 767 1 1487
2 770 1 1490
2 771 1 1490
2 773 1 1493
2 774 1 1493
2 775 1 1496
2 776 1 1496
2 777 1 1499
2 778 1 1499
2 780 1 1502
2 781 1 1502
2 783 1 1520
2 784 1 1520
2 785 1 1520
2 787 1 1562
2 788 1 1562
2 789 1 1562
2 790 1 1562
2 791 1 1562
2 792 1 1562
2 795 1 1562
2 796 1 1562
2 797 1 1562
2 799 1 1562
2 800 1 1562
2 801 1 1562
2 802 1 1562
2 804 1 1562
2 805 1 1562
2 806 1 1562
2 807 1 1667
2 808 1 1667
2 809 1 1670
2 810 1 1670
2 811 1 1715
2 812 1 1715
2 813 1 1718
2 814 1 1718
2 815 1 1722
2 816 1 1722
2 817 1 1738
2 818 1 1738
2 819 1 1738
2 822 1 1738
2 823 1 1738
2 824 1 1738
2 826 1 1738
2 827 1 1738
2 828 1 1747
2 830 1 1747
2 831 1 1747
2 833 1 1747
2 834 1 1747
2 837 1 1747
2 838 1 1747
2 840 1 1747
2 841 1 1756
2 843 1 1756
2 844 1 1756
2 846 1 1756
2 847 1 1761
2 849 1 1761
2 850 1 1803
2 852 1 1803
2 853 1 1806
2 855 1 1806
2 856 1 1809
2 857 1 1809
2 859 1 1812
2 860 1 1812
2 862 1 1815
2 863 1 1815
2 865 1 1818
2 866 1 1818
2 868 1 1821
2 869 1 1821
2 871 1 1824
2 872 1 1824
2 873 1 1824
2 875 1 1824
2 876 1 1824
2 878 1 1824
2 879 1 1824
2 881 1 1824
2 882 1 1833
2 884 1 1833
2 885 1 1833
2 887 1 1833
2 888 1 1833
2 893 1 1833
2 894 1 1833
2 897 1 1833
2 898 1 1870
2 899 1 1870
2 900 1 1875
2 901 1 1875
2 902 1 1880
2 903 1 1880
2 904 1 1885
2 905 1 1885
2 906 1 1890
2 907 1 1890
2 908 1 1895
2 909 1 1895
2 910 1 1900
2 911 1 1900
2 912 1 1905
2 918 1 1905
2 919 1 1909
2 921 1 1909
2 922 1 1913
2 924 1 1913
2 925 1 1913
2 927 1 1917
2 928 1 1917
2 930 1 1917
2 931 1 1917
2 933 1 1922
2 934 1 1922
2 936 1 1922
2 937 1 1926
2 939 1 1926
2 940 1 1926
2 942 1 1930
2 943 1 1930
2 945 1 1933
2 946 1 1933
2 948 1 1936
2 949 1 1936
2 951 1 1983
2 952 1 1983
2 954 1 2038
2 955 1 2038
2 957 1 2038
2 958 1 2038
2 960 1 2043
2 961 1 2043
2 963 1 2043
2 964 1 2043
2 966 1 2043
2 967 1 2043
2 968 1 2043
2 969 1 2043
2 970 1 2052
2 971 1 2052
2 972 1 2052
2 973 1 2052
2 974 1 2057
2 975 1 2057
2 976 1 2057
2 977 1 2057
2 978 1 2057
2 979 1 2057
2 980 1 2057
2 981 1 2057
2 982 1 2068
2 983 1 2068
2 984 1 2073
2 985 1 2073
2 986 1 2078
2 987 1 2078
2 988 1 2083
2 989 1 2083
2 990 1 2088
2 991 1 2088
2 992 1 2093
2 993 1 2093
2 994 1 2098
2 995 1 2098
2 996 1 2103
2 997 1 2103
2 998 1 2158
2 999 1 2158
2 1000 1 2158
2 1001 1 2158
2 1002 1 2158
2 1003 1 2158
2 1004 1 2158
2 1005 1 2158
2 1006 1 2158
2 1007 1 2158
2 1008 1 2158
2 1009 1 2158
2 1010 1 2158
2 1011 1 2158
2 1012 1 2158
2 1013 1 2158
2 1014 1 2175
2 1015 1 2175
2 1016 1 2185
2 1017 1 2185
2 1018 1 2188
2 1019 1 2188
2 1020 1 2191
2 1021 1 2191
2 1022 1 2194
2 1023 1 2194
2 1024 1 2197
2 1025 1 2197
2 1026 1 2200
2 1027 1 2200
2 1028 1 2203
2 1029 1 2203
2 1030 1 2206
2 1031 1 2206
2 1032 1 2212
2 1033 1 2212
2 1034 1 2212
2 1035 1 2212
2 1036 1 2212
2 1037 1 2212
2 1038 1 2212
2 1039 1 2212
2 1040 1 2221
2 1041 1 2221
2 1042 1 2221
2 1043 1 2221
2 1044 1 2221
2 1045 1 2221
2 1046 1 2221
2 1047 1 2221
2 1048 1 2270
2 1049 1 2270
2 1050 1 2277
2 1051 1 2277
2 1052 1 2282
2 1053 1 2282
2 1054 1 2287
2 1055 1 2287
2 1056 1 2294
2 1057 1 2294
2 1058 1 2299
2 1059 1 2299
2 1060 1 2304
2 1061 1 2304
2 1062 1 2307
2 1063 1 2307
2 1064 1 2310
2 1065 1 2310
2 1066 1 2313
2 1068 1 2313
2 1069 1 2316
2 1070 1 2316
2 1071 1 2319
2 1072 1 2319
2 1073 1 2322
2 1074 1 2322
2 1075 1 2325
2 1076 1 2325
2 1077 1 2328
2 1078 1 2328
2 1079 1 2331
2 1080 1 2331
2 1081 1 2334
2 1082 1 2334
2 1083 1 2376
2 1084 1 2376
2 1085 1 2379
2 1086 1 2379
2 1087 1 2471
2 1088 1 2471
2 1089 1 2483
2 1090 1 2483
2 1091 1 2488
2 1092 1 2488
2 1093 1 2488
2 1094 1 2488
2 1095 1 2488
2 1096 1 2488
2 1097 1 2488
2 1098 1 2488
2 1099 1 2497
2 1100 1 2497
2 1101 1 2497
2 1102 1 2497
2 1103 1 2497
2 1104 1 2497
2 1105 1 2497
2 1106 1 2497
2 1107 1 2506
2 1108 1 2506
2 1109 1 2506
2 1110 1 2506
2 1111 1 2506
2 1112 1 2506
2 1113 1 2506
2 1114 1 2506
2 1115 1 2515
2 1116 1 2515
2 1118 1 2515
2 1119 1 2515
2 1120 1 2515
2 1121 1 2515
2 1122 1 2515
2 1123 1 2515
2 1124 1 2524
2 1125 1 2524
2 1126 1 2524
2 1127 1 2524
2 1128 1 2524
2 1129 1 2524
2 1130 1 2524
2 1131 1 2524
2 1132 1 2533
2 1133 1 2533
2 1134 1 2533
2 1135 1 2533
2 1136 1 2533
2 1137 1 2533
2 1138 1 2533
2 1139 1 2533
2 1140 1 2542
2 1141 1 2542
2 1142 1 2542
2 1143 1 2542
2 1144 1 2542
2 1145 1 2542
2 1146 1 2542
2 1147 1 2542
2 1148 1 2551
2 1149 1 2551
2 1150 1 2551
2 1151 1 2551
2 1152 1 2551
2 1153 1 2551
2 1154 1 2551
2 1155 1 2551
2 1156 1 2560
2 1157 1 2560
2 1158 1 2560
2 1159 1 2560
2 1160 1 2560
2 1161 1 2560
2 1162 1 2560
2 1163 1 2560
2 1164 1 2569
2 1165 1 2569
2 1166 1 2569
2 1167 1 2569
2 1168 1 2569
2 1169 1 2569
2 1170 1 2569
2 1171 1 2569
2 1172 1 2578
2 1173 1 2578
2 1174 1 2578
2 1175 1 2578
2 1176 1 2578
2 1177 1 2578
2 1178 1 2578
2 1180 1 2578
2 1181 1 2587
2 1182 1 2587
2 1183 1 2587
2 1184 1 2587
2 1185 1 2587
2 1186 1 2587
2 1187 1 2587
2 1188 1 2587
2 1189 1 2596
2 1190 1 2596
2 1191 1 2596
2 1192 1 2596
2 1193 1 2596
2 1194 1 2596
2 1195 1 2596
2 1198 1 2596
2 1199 1 2605
2 1200 1 2605
2 1201 1 2605
2 1203 1 2605
2 1204 1 2605
2 1205 1 2605
2 1206 1 2605
2 1207 1 2605
2 1208 1 2614
2 1209 1 2614
2 1210 1 2614
2 1211 1 2614
2 1212 1 2614
2 1213 1 2614
2 1214 1 2614
2 1215 1 2614
2 1216 1 2623
2 1217 1 2623
2 1218 1 2623
2 1220 1 2623
2 1221 1 2623
2 1222 1 2623
2 1223 1 2623
2 1224 1 2623
2 1225 1 2648
2 1226 1 2648
2 1227 1 2648
2 1228 1 2652
2 1229 1 2652
2 1230 1 2652
2 1231 1 2656
2 1232 1 2656
2 1233 1 2659
2 1234 1 2659
2 1235 1 2662
2 1236 1 2662
2 1237 1 2662
2 1238 1 2666
2 1239 1 2666
2 1240 1 2666
2 1241 1 2670
2 1242 1 2670
2 1243 1 2673
2 1244 1 2673
2 1245 1 2673
2 1246 1 2677
2 1247 1 2677
2 1248 1 2677
2 1249 1 2681
2 1265 1 2681
2 1266 1 2684
2 1269 1 2684
2 1270 1 2684
2 1274 1 2688
2 1275 1 2688
2 1277 1 2688
2 1278 1 2692
2 1280 1 2692
2 1281 1 2692
2 1282 1 2692
2 1283 1 2697
2 1284 1 2697
2 1285 1 2697
2 1286 1 2697
2 1287 1 2702
2 1288 1 2702
2 1289 1 2702
2 1290 1 2706
2 1291 1 2706
2 1292 1 2706
2 1293 1 2710
2 1294 1 2710
2 1295 1 2710
2 1296 1 2710
2 1297 1 2715
2 1299 1 2715
2 1300 1 2715
2 1301 1 2719
2 1303 1 2719
2 1304 1 2719
2 1305 1 2723
2 1307 1 2723
2 1308 1 2723
2 1309 1 2723
2 1310 1 2758
2 1311 1 2758
2 1312 1 2761
2 1313 1 2761
2 1314 1 2764
2 1316 1 2764
2 1317 1 2967
2 1318 1 2967
2 1319 1 2970
2 1320 1 2970
2 1321 1 2973
2 1323 1 2973
2 1324 1 2973
2 1326 1 2977
2 1327 1 2977
2 1329 1 3112
2 1330 1 3112
2 1332 1 3115
2 1333 1 3115
2 1335 1 3119
2 1336 1 3119
2 1341 1 3122
2 1342 1 3122
2 1354 1 3125
2 1355 1 3125
2 1356 1 3128
2 1357 1 3128
2 1359 1 3131
2 1360 1 3131
2 1361 1 3135
2 1362 1 3135
2 1364 1 3138
2 1365 1 3138
2 1367 1 3142
2 1368 1 3142
2 1370 1 3145
2 1371 1 3145
2 1372 1 3149
2 1373 1 3149
2 1374 1 3152
2 1375 1 3152
2 1376 1 3155
2 1377 1 3155
2 1378 1 3158
2 1379 1 3158
2 1380 1 3161
2 1381 1 3161
2 1382 1 3165
2 1383 1 3165
2 1385 1 3168
2 1386 1 3168
2 1387 1 3172
2 1388 1 3172
2 1389 1 3175
2 1390 1 3175
2 1391 1 3178
2 1392 1 3178
2 1393 1 3181
2 1394 1 3181
2 1395 1 3184
2 1396 1 3184
2 1397 1 3187
2 1398 1 3187
2 1399 1 3384
2 1400 1 3384
2 1410 1 3407
2 1411 1 3407
2 1412 1 3410
2 1413 1 3410
2 1414 1 3415
2 1415 1 3415
2 1416 1 3415
2 1417 1 3419
2 1418 1 3419
2 1419 1 3419
2 1420 1 3423
2 1421 1 3423
2 1422 1 3426
2 1423 1 3426
2 1424 1 3431
2 1425 1 3431
2 1428 1 3434
2 1429 1 3434
2 1430 1 3439
2 1431 1 3439
2 1432 1 3442
2 1433 1 3442
2 1434 1 3447
2 1435 1 3447
2 1436 1 3447
2 1437 1 3451
2 1438 1 3451
2 1439 1 3451
2 1440 1 3455
2 1441 1 3455
2 1442 1 3458
2 1443 1 3458
2 1444 1 3463
2 1445 1 3463
2 1446 1 3466
2 1447 1 3466
2 1448 1 3472
2 1449 1 3472
2 1450 1 3475
2 1451 1 3475
2 1453 1 3478
2 1454 1 3478
2 1455 1 3481
2 1456 1 3481
2 1457 1 3484
2 1458 1 3484
2 1462 1 3487
2 1463 1 3487
2 1465 1 3490
2 1466 1 3490
2 1472 1 3493
2 1473 1 3493
2 1476 1 3496
2 1477 1 3496
2 1479 1 3499
2 1480 1 3499
2 1482 1 3502
2 1483 1 3502
2 1485 1 3505
2 1486 1 3505
2 1488 1 3508
2 1489 1 3508
2 1491 1 3511
2 1492 1 3511
2 1494 1 3514
2 1495 1 3514
2 1497 1 3517
2 1498 1 3517
2 1500 1 3520
2 1501 1 3520
2 1503 1 3523
2 1504 1 3523
2 1506 1 3645
2 1513 1 3645
2 1514 1 3648
2 1515 1 3648
2 1516 1 3654
2 1517 1 3654
2 1518 1 3658
2 1519 1 3658
2 1521 1 3664
2 1522 1 3664
2 1523 1 3667
2 1524 1 3667
2 1525 1 3673
2 1526 1 3673
2 1527 1 3677
2 1528 1 3677
2 1529 1 3682
2 1530 1 3682
2 1531 1 3690
2 1532 1 3690
2 1533 1 3697
2 1534 1 3697
2 1535 1 3700
2 1536 1 3700
2 1537 1 3721
2 1538 1 3721
2 1539 1 3721
2 1540 1 3721
2 1541 1 3721
2 1542 1 3734
2 1543 1 3734
2 1544 1 3734
2 1545 1 3740
2 1546 1 3740
2 1547 1 3743
2 1548 1 3743
2 1549 1 3743
2 1550 1 3743
2 1551 1 3743
2 1552 1 3756
2 1553 1 3756
2 1554 1 3756
2 1555 1 3762
2 1556 1 3762
2 1557 1 3786
2 1558 1 3786
2 1559 1 3800
2 1560 1 3800
2 1561 1 3809
2 1563 1 3809
2 1564 1 3812
2 1565 1 3812
2 1566 1 3815
2 1567 1 3815
2 1568 1 3818
2 1569 1 3818
2 1570 1 3821
2 1571 1 3821
2 1572 1 3824
2 1573 1 3824
2 1574 1 3827
2 1575 1 3827
2 1576 1 3830
2 1577 1 3830
2 1578 1 3838
2 1601 1 3838
2 1602 1 3838
2 1603 1 3838
2 1604 1 3845
2 1605 1 3845
2 1606 1 3845
2 1607 1 3845
2 1608 1 3850
2 1609 1 3850
2 1610 1 3855
2 1611 1 3855
2 1612 1 3858
2 1613 1 3858
2 1614 1 3861
2 1615 1 3861
2 1616 1 3865
2 1617 1 3865
2 1618 1 3868
2 1619 1 3868
2 1620 1 3913
2 1621 1 3913
2 1622 1 3917
2 1623 1 3917
2 1624 1 3921
2 1625 1 3921
2 1626 1 3926
2 1627 1 3926
2 1628 1 3926
2 1629 1 3932
2 1630 1 3932
2 1631 1 3937
2 1632 1 3937
2 1633 1 3940
2 1634 1 3940
2 1635 1 3950
2 1636 1 3950
2 1637 1 3953
2 1638 1 3953
2 1639 1 3956
2 1640 1 3956
2 1641 1 3959
2 1642 1 3959
2 1651 1 3962
2 1652 1 3962
2 1653 1 3965
2 1654 1 3965
2 1655 1 3968
2 1656 1 3968
2 1657 1 3971
2 1658 1 3971
2 1659 1 3974
2 1660 1 3974
2 1661 1 3977
2 1662 1 3977
2 1663 1 3980
2 1664 1 3980
2 1665 1 3983
2 1666 1 3983
2 1668 1 3992
2 1669 1 3992
2 1671 1 3996
2 1672 1 3996
2 1681 1 4035
2 1682 1 4035
2 1683 1 4059
2 1684 1 4059
2 1685 1 4062
2 1686 1 4062
2 1687 1 4067
2 1688 1 4067
2 1689 1 4070
2 1690 1 4070
2 1695 1 4091
2 1696 1 4091
2 1697 1 4094
2 1698 1 4094
2 1699 1 4094
2 1700 1 4116
2 1701 1 4116
2 1702 1 4119
2 1703 1 4119
2 1704 1 4123
2 1705 1 4123
2 1706 1 4128
2 1707 1 4128
2 1708 1 4128
2 1709 1 4128
2 1710 1 4128
2 1711 1 4139
2 1712 1 4139
2 1716 1 4142
2 1717 1 4142
2 1719 1 4167
2 1720 1 4167
2 1723 1 4167
2 1724 1 4167
2 1732 1 4167
2 1733 1 4167
2 1734 1 4174
2 1739 1 4174
2 1740 1 4174
2 1741 1 4174
2 1742 1 4182
2 1743 1 4182
2 1744 1 4186
2 1745 1 4186
2 1746 1 4197
2 1748 1 4197
2 1749 1 4200
2 1750 1 4200
2 1751 1 4203
2 1752 1 4203
2 1753 1 4203
2 1754 1 4203
2 1755 1 4203
2 1757 1 4209
2 1758 1 4209
2 1759 1 4209
2 1760 1 4213
2 1762 1 4213
2 1763 1 4213
2 1771 1 4213
2 1772 1 4218
2 1773 1 4218
2 1774 1 4218
2 1775 1 4218
2 1776 1 4223
2 1777 1 4223
2 1778 1 4223
2 1779 1 4223
2 1780 1 4242
2 1781 1 4242
2 1782 1 4247
2 1783 1 4247
2 1784 1 4284
2 1785 1 4284
2 1786 1 4287
2 1804 1 4287
2 1805 1 4287
2 1807 1 4296
2 1808 1 4296
2 1810 1 4305
2 1811 1 4305
2 1813 1 4305
2 1814 1 4305
2 1816 1 4310
2 1817 1 4310
2 1819 1 4310
2 1820 1 4319
2 1822 1 4319
2 1823 1 4331
2 1825 1 4331
2 1826 1 4335
2 1827 1 4335
2 1828 1 4338
2 1829 1 4338
2 1830 1 4341
2 1831 1 4341
2 1832 1 4344
2 1834 1 4344
2 1835 1 4347
2 1836 1 4347
2 1837 1 4350
2 1838 1 4350
2 1839 1 4353
2 1840 1 4353
2 1841 1 4356
2 1865 1 4356
2 1866 1 4359
2 1867 1 4359
2 1868 1 4362
2 1871 1 4362
2 1872 1 4365
2 1876 1 4365
2 1877 1 4368
2 1881 1 4368
2 1882 1 4371
2 1886 1 4371
2 1887 1 4387
2 1891 1 4387
2 1892 1 4390
2 1896 1 4390
2 1897 1 4398
2 1901 1 4398
2 1902 1 4413
2 1906 1 4413
2 1907 1 4416
2 1910 1 4416
2 1911 1 4421
2 1914 1 4421
2 1915 1 4427
2 1916 1 4427
2 1918 1 4430
2 1919 1 4430
2 1920 1 4435
2 1921 1 4435
2 1923 1 4443
2 1924 1 4443
2 1925 1 4458
2 1927 1 4458
2 1928 1 4465
2 1929 1 4465
2 1931 1 4468
2 1932 1 4468
2 1934 1 4472
2 1935 1 4472
2 1937 1 4475
2 1938 1 4475
2 1948 1 4479
2 1949 1 4479
2 1950 1 4493
2 1951 1 4493
2 1952 1 4498
2 1953 1 4498
2 1954 1 4503
2 1955 1 4503
2 1956 1 4531
2 1957 1 4531
2 1958 1 4534
2 1959 1 4534
2 1962 1 4537
2 1963 1 4537
2 1964 1 4540
2 1965 1 4540
2 1967 1 4549
2 1968 1 4549
2 1969 1 4559
2 1970 1 4559
2 1971 1 4564
2 1972 1 4564
2 1973 1 4564
2 1974 1 4569
2 1975 1 4569
2 1976 1 4576
2 1977 1 4576
2 1978 1 4581
2 1979 1 4581
2 1980 1 4584
2 1984 1 4584
2 1985 1 4593
2 1992 1 4593
2 1993 1 4599
2 1994 1 4599
2 1995 1 4613
2 1996 1 4613
2 1997 1 4616
2 1998 1 4616
2 1999 1 4619
2 2000 1 4619
2 2001 1 4623
2 2002 1 4623
2 2003 1 4644
2 2004 1 4644
2 2005 1 4647
2 2006 1 4647
2 2007 1 4650
2 2008 1 4650
2 2009 1 4656
2 2010 1 4656
2 2011 1 4659
2 2012 1 4659
2 2013 1 4664
2 2014 1 4664
2 2015 1 4691
2 2016 1 4691
2 2017 1 4694
2 2018 1 4694
2 2019 1 4697
2 2020 1 4697
2 2021 1 4700
2 2039 1 4700
2 2040 1 4711
2 2041 1 4711
2 2042 1 4717
2 2044 1 4717
2 2045 1 4717
2 2046 1 4722
2 2047 1 4722
2 2048 1 4722
2 2049 1 4727
2 2050 1 4727
2 2051 1 4730
2 2053 1 4730
2 2054 1 4740
2 2055 1 4740
2 2056 1 4743
2 2058 1 4743
2 2059 1 4743
2 2060 1 4757
2 2061 1 4757
2 2062 1 4757
2 2063 1 4769
2 2064 1 4769
2 2065 1 4772
2 2066 1 4772
2 2067 1 4775
2 2069 1 4775
2 2070 1 4794
2 2071 1 4794
2 2072 1 4797
2 2074 1 4797
2 2075 1 4800
2 2076 1 4800
2 2077 1 4805
2 2079 1 4805
2 2080 1 4808
2 2081 1 4808
2 2082 1 4812
2 2084 1 4812
2 2085 1 4818
2 2086 1 4818
2 2087 1 4818
2 2089 1 4823
2 2090 1 4823
2 2091 1 4831
2 2092 1 4831
2 2094 1 4838
2 2095 1 4838
2 2096 1 4844
2 2097 1 4844
2 2099 1 4847
2 2100 1 4847
2 2101 1 4850
2 2102 1 4850
2 2104 1 4854
2 2105 1 4854
2 2106 1 4876
2 2107 1 4876
2 2108 1 4876
2 2109 1 4880
2 2110 1 4880
2 2111 1 4889
2 2112 1 4889
2 2113 1 4907
2 2114 1 4907
2 2115 1 4913
2 2116 1 4913
2 2117 1 4916
2 2118 1 4916
2 2119 1 4921
2 2120 1 4921
2 2129 1 4937
2 2130 1 4937
2 2131 1 4940
2 2132 1 4940
2 2140 1 4946
2 2159 1 4946
2 2160 1 4954
2 2161 1 4954
2 2162 1 4957
2 2163 1 4957
2 2164 1 4973
2 2165 1 4973
2 2166 1 4985
2 2167 1 4985
2 2168 1 4988
2 2169 1 4988
2 2170 1 4991
2 2171 1 4991
2 2172 1 4996
2 2173 1 4996
2 2174 1 4999
2 2176 1 4999
2 2177 1 5010
2 2182 1 5010
2 2186 1 5013
2 2187 1 5013
2 2189 1 5018
2 2190 1 5018
2 2192 1 5021
2 2193 1 5021
2 2195 1 5030
2 2196 1 5030
2 2198 1 5039
2 2199 1 5039
2 2201 1 5042
2 2202 1 5042
2 2204 1 5050
2 2205 1 5050
2 2207 1 5050
2 2208 1 5050
2 2213 1 5055
2 2214 1 5055
2 2215 1 5058
2 2216 1 5058
2 2217 1 5061
2 2218 1 5061
2 2219 1 5066
2 2220 1 5066
2 2222 1 5070
2 2223 1 5070
2 2224 1 5080
2 2225 1 5080
2 2226 1 5080
2 2227 1 5080
2 2228 1 5085
2 2229 1 5085
2 2246 1 5111
2 2247 1 5111
2 2248 1 5114
2 2249 1 5114
2 2250 1 5117
2 2251 1 5117
2 2252 1 5122
2 2253 1 5122
2 2254 1 5128
2 2255 1 5128
2 2256 1 5133
2 2257 1 5133
2 2258 1 5139
2 2259 1 5139
2 2260 1 5145
2 2261 1 5145
2 2262 1 5151
2 2263 1 5151
2 2264 1 5154
2 2265 1 5154
2 2266 1 5160
2 2267 1 5160
2 2268 1 5163
2 2269 1 5163
2 2271 1 5174
2 2272 1 5174
2 2273 1 5177
2 2274 1 5177
2 2275 1 5184
2 2276 1 5184
2 2278 1 5188
2 2279 1 5188
2 2280 1 5205
2 2281 1 5205
2 2283 1 5209
2 2284 1 5209
2 2285 1 5228
2 2286 1 5228
2 2288 1 5236
2 2289 1 5236
2 2290 1 5236
2 2291 1 5250
2 2292 1 5250
2 2293 1 5254
2 2295 1 5254
2 2296 1 5258
2 2297 1 5258
2 2298 1 5266
2 2300 1 5266
2 2301 1 5269
2 2302 1 5269
2 2303 1 5279
2 2305 1 5279
2 2306 1 5289
2 2308 1 5289
2 2309 1 5292
2 2311 1 5292
2 2312 1 5298
2 2314 1 5298
2 2315 1 5303
2 2317 1 5303
2 2318 1 5306
2 2320 1 5306
2 2321 1 5309
2 2323 1 5309
2 2324 1 5324
2 2326 1 5324
2 2327 1 5327
2 2329 1 5327
2 2330 1 5332
2 2332 1 5332
2 2333 1 5335
2 2335 1 5335
