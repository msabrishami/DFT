1	1	0	18	0	
1	13	0	9	0	
1	20	0	15	0	
1	33	0	22	0	
1	41	0	3	0	
1	45	0	5	0	
1	50	0	16	0	
1	58	0	19	0	
1	68	0	20	0	
1	77	0	17	0	
1	87	0	17	0	
1	97	0	19	0	
1	107	0	18	0	
1	116	0	15	0	
1	124	0	1	0	
1	125	0	2	0	
1	128	0	3	0	
1	132	0	4	0	
1	137	0	5	0	
1	143	0	6	0	
1	150	0	8	0	
1	159	0	9	0	
1	169	0	9	0	
1	179	0	11	0	
1	190	0	10	0	
1	200	0	12	0	
1	213	0	8	0	
1	222	0	1	0	
1	223	0	2	0	
1	226	0	6	0	
1	232	0	6	0	
1	238	0	6	0	
1	244	0	6	0	
1	250	0	7	0	
1	257	0	7	0	
1	264	0	6	0	
1	270	0	4	0	
1	274	0	8	0	
1	283	0	10	0	
1	294	0	8	0	
1	303	0	7	0	
1	311	0	5	0	
1	317	0	4	0	
1	322	0	3	0	
1	326	0	2	0	
1	329	0	1	0	
1	330	0	13	0	
1	343	0	6	0	
1	349	0	1	0	
1	350	0	2	0	
0	665	5	5	1	5434	
0	679	5	4	1	5450	
0	686	5	4	1	5469	
0	702	5	4	1	5489	
0	724	5	3	1	5506	
0	736	5	4	1	5523	
0	749	5	4	1	5542	
0	763	5	5	1	5560	
0	768	3	1	2	5695	5702	
0	769	5	2	1	5362	
0	779	5	2	1	5363	
0	786	5	6	1	5380	
0	793	7	1	2	5381	5389	
0	794	5	3	1	5390	
0	803	5	16	1	5391	
0	820	5	1	1	5404	
0	825	5	20	1	5405	
0	829	7	2	2	5406	5426	
0	832	5	4	1	5427	
0	835	3	1	2	5428	5429	
0	839	5	4	1	5430	
0	842	5	2	1	5435	
0	848	5	2	1	5451	
0	854	5	3	1	5470	
0	861	5	2	1	5507	
0	867	5	2	1	5524	
0	870	5	3	1	5543	
0	883	5	2	1	5392	
0	889	5	1	1	5642	
0	890	7	1	2	5393	5643	
0	891	6	1	2	5394	5644	
0	892	7	3	2	5395	5621	
0	895	5	1	1	5396	
0	896	3	16	2	349	5407	
0	913	6	1	2	5364	5382	
0	914	6	1	3	5365	5397	5408	
0	915	5	1	1	5398	
0	916	5	1	1	5409	
0	920	5	2	1	5654	
0	1067	7	1	2	5688	768	
0	1117	3	16	2	820	5399	
0	1179	3	1	2	895	5612	
0	1196	5	1	1	793	
0	1197	3	4	2	915	5366	
0	1202	7	16	2	913	914	
0	1219	3	4	2	916	5367	
0	1250	7	1	3	5872	5874	5876	
0	1251	6	1	2	5664	5436	
0	1252	6	1	2	5670	5452	
0	1253	6	1	2	5676	5471	
0	1254	6	1	2	5682	5490	
0	1255	6	1	2	5689	5508	
0	1256	6	1	2	5696	5525	
0	1257	6	1	2	5703	5544	
0	1258	6	1	2	5708	5561	
0	1259	5	1	1	5665	
0	1260	5	1	1	5671	
0	1261	5	1	1	5677	
0	1262	5	1	1	5683	
0	1263	6	1	2	5785	5789	
0	1264	6	2	2	5800	5804	
0	1267	6	1	2	5472	5491	
0	1271	5	1	1	5453	
0	1272	5	1	1	5526	
0	1306	7	8	2	5815	835	
0	1315	7	6	3	5816	5431	5864	
0	1322	7	2	2	5813	5432	
0	1325	7	2	3	5368	5817	5400	
0	1328	6	2	3	5369	5818	5401	
0	1331	6	2	2	5370	5819	
0	1337	6	1	3	5383	5823	5433	
0	1338	6	1	3	5873	5875	5877	
0	1339	5	1	1	5454	
0	1340	7	2	3	5879	5881	5883	
0	1343	6	1	3	5880	5882	5884	
0	1344	5	1	1	5527	
0	1345	5	1	1	5826	
0	1346	5	1	1	5827	
0	1347	5	1	1	5828	
0	1348	5	1	1	5829	
0	1349	5	1	1	5830	
0	1350	5	1	1	5831	
0	1351	5	1	1	5832	
0	1352	5	1	1	5833	
0	1353	3	4	2	5886	5632	
0	1358	4	4	2	5887	5633	
0	1366	5	2	1	5888	
0	1401	5	1	1	5891	
0	1402	5	1	1	5892	
0	1403	5	1	1	5893	
0	1404	5	1	1	5894	
0	1405	5	1	1	5895	
0	1406	5	1	1	5896	
0	1407	5	1	1	5897	
0	1408	5	1	1	5898	
0	1409	3	16	2	5371	1196	
0	1426	5	1	1	5862	
0	1427	5	1	1	5863	
0	1452	7	6	3	5814	5384	5824	
0	1459	5	1	1	5622	
0	1460	5	1	1	5759	
0	1461	3	2	2	5907	5772	
0	1464	4	3	2	5908	5773	
0	1467	5	1	1	5690	
0	1468	5	1	1	5697	
0	1469	5	1	1	5704	
0	1470	5	1	1	5709	
0	1474	5	1	1	5437	
0	1505	6	1	2	5793	1250	
0	1507	7	1	4	1251	1252	1253	1254	
0	1508	7	1	4	1255	1256	1257	1258	
0	1509	6	1	2	5672	1259	
0	1510	6	1	2	5666	1260	
0	1511	6	1	2	5684	1261	
0	1512	6	1	2	5678	1262	
0	1520	7	3	2	5438	1263	
0	1562	7	16	2	5372	1337	
0	1579	5	1	1	5909	
0	1580	7	1	2	5834	5910	
0	1581	7	1	2	1338	1345	
0	1582	5	1	1	5911	
0	1583	7	1	2	5835	5912	
0	1584	5	1	1	5913	
0	1585	7	1	2	5836	5914	
0	1586	7	1	2	5878	1347	
0	1587	5	1	1	5915	
0	1588	7	1	2	5837	5916	
0	1589	7	1	2	5492	1348	
0	1590	5	1	1	5917	
0	1591	7	1	2	5838	5918	
0	1592	7	1	2	1343	1349	
0	1593	5	1	1	5919	
0	1594	7	1	2	5839	5920	
0	1595	5	1	1	5921	
0	1596	7	1	2	5840	5922	
0	1597	7	1	2	5885	1351	
0	1598	5	1	1	5923	
0	1599	7	1	2	5841	5924	
0	1600	7	1	2	5562	1352	
0	1643	7	1	2	222	1401	
0	1644	7	1	2	5662	1402	
0	1645	7	1	2	5667	1403	
0	1646	7	1	2	5673	1404	
0	1647	7	1	2	5679	1405	
0	1648	7	1	2	5685	1406	
0	1649	7	1	2	5691	1407	
0	1650	7	1	2	5698	1408	
0	1667	7	5	3	5373	5385	1426	
0	1670	7	5	3	5374	5386	1427	
0	1673	5	1	1	5929	
0	1674	5	1	1	5930	
0	1675	5	1	1	5931	
0	1676	5	1	1	5932	
0	1677	5	1	1	5933	
0	1678	5	1	1	5934	
0	1679	5	1	1	5935	
0	1680	5	1	1	5936	
0	1691	6	1	2	5699	1467	
0	1692	6	1	2	5692	1468	
0	1693	6	1	2	5710	1469	
0	1694	6	1	2	5705	1470	
3	1713	5	0	1	1505	
0	1714	7	1	2	5509	5949	
0	1715	6	4	2	1509	1510	
0	1718	6	4	2	1511	1512	
0	1721	6	1	2	1507	1508	
0	1722	7	2	2	5808	5973	
0	1725	6	1	2	5809	5974	
0	1726	5	1	1	5780	
0	1727	6	1	2	5473	1271	
0	1728	5	1	1	5474	
0	1729	7	1	2	5475	5781	
0	1730	6	1	2	5545	1272	
0	1731	5	1	1	5546	
0	1735	6	1	2	5510	5950	
0	1736	5	1	1	5868	
0	1737	5	1	1	5869	
0	1738	6	8	2	5967	5410	
0	1747	6	8	2	5968	5842	
0	1756	6	4	3	5375	5387	5402	
0	1761	6	18	4	5376	5820	5403	5865	
0	1764	6	1	2	5476	1339	
0	1765	5	1	1	5477	
0	1766	6	1	2	5547	1344	
0	1767	5	1	1	5548	
0	1768	5	1	1	5969	
0	1769	5	1	1	5377	
0	1770	5	1	1	5971	
0	1787	7	1	2	5455	1579	
0	1788	7	1	2	5595	1580	
0	1789	7	1	2	5478	1582	
0	1790	7	1	2	5603	1583	
0	1791	7	1	2	5493	1584	
0	1792	7	1	2	5439	1585	
0	1793	7	1	2	5511	1587	
0	1794	7	1	2	5456	1588	
0	1795	7	1	2	5528	1590	
0	1796	7	1	2	5479	1591	
0	1797	7	1	2	5549	1593	
0	1798	7	1	2	5494	1594	
0	1799	7	1	2	5563	1595	
0	1800	7	1	2	5512	1596	
0	1801	7	1	2	5720	1598	
0	1802	7	1	2	5529	1599	
0	1803	7	2	2	5645	5889	
0	1806	7	2	2	889	5890	
0	1809	7	2	2	890	5983	
0	1812	7	2	2	891	5984	
0	1815	6	2	2	5843	5866	
0	1818	6	2	2	5411	5867	
0	1821	6	16	3	5378	5388	1179	
0	1824	6	8	3	5821	5825	5844	
0	1833	6	8	2	5822	5845	
0	1842	5	1	1	5412	
0	1843	5	1	1	5413	
0	1844	5	1	1	5414	
0	1845	5	1	1	5415	
0	1846	5	1	1	5416	
0	1847	5	1	1	5417	
0	1848	5	1	1	5418	
0	1849	5	1	1	5846	
0	1850	7	1	2	5847	5899	
0	1851	5	1	1	5848	
0	1852	7	1	2	5849	5900	
0	1853	5	1	1	5850	
0	1854	7	1	2	5851	5901	
0	1855	5	1	1	5852	
0	1856	7	1	2	5853	5902	
0	1857	5	1	1	5854	
0	1858	7	1	2	5855	5903	
0	1859	5	1	1	5856	
0	1860	7	1	2	5857	5904	
0	1861	5	1	1	5858	
0	1862	7	1	2	5859	5905	
0	1863	5	1	1	5860	
0	1864	7	1	2	5861	5906	
0	1869	7	1	2	5937	5985	
0	1870	4	2	2	5440	5986	
0	1873	5	1	1	5951	
0	1874	7	1	2	5938	5987	
0	1875	4	2	2	5457	5988	
0	1878	5	1	1	5952	
0	1879	7	1	2	5939	5989	
0	1880	4	2	2	5480	5990	
0	1883	5	1	1	5953	
0	1884	7	1	2	5940	5991	
0	1885	4	2	2	5495	5992	
0	1888	5	1	1	5954	
0	1889	7	1	2	5941	5993	
0	1890	4	2	2	5513	5994	
0	1893	5	1	1	5965	
0	1894	7	1	2	5942	5995	
0	1895	4	2	2	5530	5996	
0	1898	5	1	1	5959	
0	1899	7	1	2	5943	5997	
0	1900	4	2	2	5550	5998	
0	1903	5	1	1	5960	
0	1904	7	1	2	5944	5999	
0	1905	4	2	2	5564	6000	
0	1908	5	1	1	5961	
0	1909	7	2	2	6001	5655	
0	1912	6	1	2	6002	5656	
0	1913	7	3	3	6003	5657	5774	
0	1917	6	5	3	6004	5658	5775	
0	1922	7	3	3	6005	5659	5776	
0	1926	6	3	3	6006	5660	5777	
0	1933	6	2	2	1691	1692	
0	1936	6	2	2	1693	1694	
0	1939	5	1	1	5786	
0	1940	6	1	2	5787	1474	
0	1941	5	1	1	5790	
0	1942	5	1	1	5794	
0	1943	5	1	1	5797	
0	1944	5	1	1	5801	
0	1945	5	1	1	5805	
0	1946	5	1	1	5810	
3	1947	5	0	1	1714	
0	1960	6	1	2	5458	1728	
0	1961	6	1	2	5531	1731	
0	1966	7	1	2	6012	5870	
0	1981	6	1	2	5459	1765	
0	1982	6	1	2	5532	1767	
0	1983	7	2	2	1067	1768	
0	1986	3	1	3	1581	1787	1788	
0	1987	3	1	3	1586	1791	1792	
0	1988	3	1	3	1589	1793	1794	
0	1989	3	1	3	1592	1795	1796	
0	1990	3	1	3	1597	1799	1800	
0	1991	3	1	3	1600	1801	1802	
0	2022	7	1	2	5496	1849	
0	2023	7	1	2	5663	1850	
0	2024	7	1	2	5514	1851	
0	2025	7	1	2	5668	1852	
0	2026	7	1	2	5533	1853	
0	2027	7	1	2	5674	1854	
0	2028	7	1	2	5551	1855	
0	2029	7	1	2	5680	1856	
0	2030	7	1	2	5565	1857	
0	2031	7	1	2	5686	1858	
0	2032	7	1	2	5721	1859	
0	2033	7	1	2	5693	1860	
0	2034	7	1	2	5730	1861	
0	2035	7	1	2	5700	1862	
0	2036	7	1	2	5738	1863	
0	2037	7	1	2	5706	1864	
0	2043	5	8	1	6031	
0	2057	5	8	1	6036	
0	2068	7	2	3	5441	5925	1869	
0	2073	7	2	3	5460	5926	1874	
0	2078	7	2	3	5481	5927	1879	
0	2083	7	2	3	5497	5928	1884	
0	2088	7	2	3	5515	5945	1889	
0	2093	7	2	3	5534	5946	1894	
0	2098	7	2	3	5552	5947	1899	
0	2103	7	2	3	5566	5948	1904	
0	2121	5	1	1	6015	
0	2122	5	1	1	6016	
0	2123	5	1	1	6017	
0	2124	5	1	1	6018	
0	2125	5	1	1	6019	
0	2126	5	1	1	6020	
0	2127	5	1	1	6021	
0	2128	5	1	1	6022	
0	2133	6	1	2	5442	1939	
0	2134	6	1	2	5795	1941	
0	2135	6	1	2	5791	1942	
0	2136	6	1	2	5802	1943	
0	2137	6	1	2	5798	1944	
0	2138	6	1	2	5811	1945	
0	2139	6	1	2	5806	1946	
0	2141	5	1	1	6165	
0	2142	5	1	1	6167	
0	2143	5	1	1	6051	
0	2144	7	1	2	6052	6059	
0	2145	5	1	1	6060	
0	2146	6	1	2	1727	1960	
0	2147	6	1	2	1730	1961	
0	2148	7	1	4	6049	1267	5782	5461	
0	2149	5	1	1	6053	
0	2150	7	1	2	6054	6061	
0	2151	5	1	1	6062	
0	2152	5	1	1	6055	
0	2153	5	1	1	6063	
0	2154	7	1	2	6056	6064	
0	2155	5	1	1	6057	
0	2156	5	1	1	6065	
0	2157	7	1	2	6058	6066	
0	2178	6	1	2	1764	1981	
0	2179	6	1	2	1766	1982	
0	2180	5	1	1	6067	
0	2181	7	1	2	6068	5970	
0	2183	5	1	1	6069	
0	2184	7	1	2	5972	6070	
0	2185	6	16	2	5979	6095	
0	2188	6	16	2	5980	6093	
0	2191	6	16	2	5975	6096	
0	2194	6	16	2	5976	6094	
0	2197	6	16	2	5981	6091	
0	2200	6	16	2	5982	6089	
0	2203	6	16	2	5977	6092	
0	2206	6	16	2	5978	6090	
0	2209	5	1	1	6097	
0	2210	5	1	1	6099	
0	2211	7	1	2	6098	6100	
0	2230	5	1	1	6125	
0	2231	5	1	1	6126	
0	2232	5	1	1	6127	
0	2233	5	1	1	6128	
0	2234	5	1	1	6117	
0	2235	5	1	1	6118	
0	2236	5	1	1	6119	
0	2237	5	1	1	6120	
0	2238	3	1	3	2022	1643	2023	
0	2239	3	1	3	2024	1644	2025	
0	2240	3	1	3	2026	1645	2027	
0	2241	3	1	3	2028	1646	2029	
0	2242	3	1	3	2030	1647	2031	
0	2243	3	1	3	2032	1648	2033	
0	2244	3	1	3	2034	1649	2035	
0	2245	3	1	3	2036	1650	2037	
0	2270	7	2	2	1986	1673	
0	2277	7	2	2	1987	1675	
0	2282	7	2	2	1988	1676	
0	2287	7	2	2	1989	1677	
0	2294	7	2	2	1990	1679	
0	2299	7	2	2	1991	1680	
0	2307	7	2	2	6009	5778	
0	2310	6	2	2	6010	5779	
0	2325	6	2	2	1940	2133	
0	2328	6	2	2	2134	2135	
0	2331	6	2	2	2136	2137	
0	2334	6	2	2	2138	2139	
0	2341	6	1	2	6168	2141	
0	2342	6	1	2	6166	2142	
0	2347	7	1	2	5799	2144	
0	2348	7	1	3	2146	5498	1726	
0	2349	7	1	2	5567	2147	
0	2350	7	1	2	2148	5871	
0	2351	7	1	2	5803	2150	
0	2352	7	1	2	1735	2153	
0	2353	7	1	2	5812	2154	
0	2354	7	1	2	1725	2156	
0	2355	7	1	2	5807	2157	
0	2374	5	1	1	2178	
0	2375	5	1	1	2179	
0	2376	7	2	2	6013	2180	
0	2379	7	2	2	1721	2181	
0	2398	7	1	2	5783	2211	
0	2417	7	1	3	6179	5669	1873	
0	2418	7	1	3	6180	5712	5955	
0	2419	7	1	2	6037	2238	
0	2420	7	1	3	6181	5675	1878	
0	2421	7	1	3	6182	5713	5956	
0	2422	7	1	2	6038	2239	
0	2425	7	1	3	6183	5681	1883	
0	2426	7	1	3	6184	5714	5957	
0	2427	7	1	2	6039	2240	
0	2430	7	1	3	6185	5687	1888	
0	2431	7	1	3	6186	5715	5958	
0	2432	7	1	2	6040	2241	
0	2435	7	1	3	6171	5694	1893	
0	2436	7	1	3	6172	5716	5966	
0	2437	7	1	2	6032	2242	
0	2438	7	1	3	6173	5701	1898	
0	2439	7	1	3	6174	5717	5962	
0	2440	7	1	2	6033	2243	
0	2443	7	1	3	6175	5707	1903	
0	2444	7	1	3	6176	5718	5963	
0	2445	7	1	2	6034	2244	
0	2448	7	1	3	6177	5711	1908	
0	2449	7	1	3	6178	5719	5964	
0	2450	7	1	2	6035	2245	
0	2467	5	1	1	6041	
0	2468	5	1	1	6045	
0	2469	5	1	1	6042	
0	2470	5	1	1	6046	
0	2471	6	5	2	2341	2342	
0	2474	5	1	1	6347	
0	2475	5	1	1	6349	
0	2476	5	1	1	6351	
0	2477	5	1	1	6353	
0	2478	3	1	2	2348	1729	
0	2481	5	1	1	6071	
0	2482	7	1	2	6072	5379	
0	2483	7	2	2	2349	2183	
0	2486	7	1	2	2374	1346	
0	2487	7	1	2	2375	1350	
0	2632	5	1	1	6101	
0	2633	7	1	2	6102	6129	
0	2634	5	1	1	6103	
0	2635	7	1	2	6104	6130	
0	2636	5	1	1	6105	
0	2637	7	1	2	6106	6131	
0	2638	5	1	1	6107	
0	2639	7	1	2	6108	6132	
0	2640	5	1	1	6109	
0	2641	7	1	2	6110	6121	
0	2642	5	1	1	6111	
0	2643	7	1	2	6112	6122	
0	2644	5	1	1	6113	
0	2645	7	1	2	6114	6123	
0	2646	5	1	1	6115	
0	2647	7	1	2	6116	6124	
0	2648	3	3	3	6331	6133	6187	
0	2652	4	3	3	6332	6134	6188	
0	2656	3	3	3	2417	2418	2419	
0	2659	3	3	3	2420	2421	2422	
0	2662	3	3	3	6333	6137	6191	
0	2666	4	3	3	6334	6138	6192	
0	2670	3	3	3	2425	2426	2427	
0	2673	3	3	3	6335	6139	6193	
0	2677	4	3	3	6336	6140	6194	
0	2681	3	3	3	2430	2431	2432	
0	2684	3	3	3	6337	6141	6195	
0	2688	4	3	3	6338	6142	6196	
0	2692	3	5	3	2435	2436	2437	
0	2697	3	5	3	2438	2439	2440	
0	2702	3	3	3	6339	6145	6199	
0	2706	4	3	3	6340	6146	6200	
0	2710	3	5	3	2443	2444	2445	
0	2715	3	3	3	6341	6147	6201	
0	2719	4	3	3	6342	6148	6202	
0	2723	3	5	3	2448	2449	2450	
0	2728	5	1	1	6154	
0	2729	5	1	1	6073	
0	2730	7	1	2	6023	6074	
0	2731	5	1	1	6075	
0	2732	7	1	2	6024	6076	
0	2733	5	1	1	6077	
0	2734	7	1	2	6025	6078	
0	2735	5	1	1	6079	
0	2736	7	1	2	6026	6080	
0	2737	5	1	1	6081	
0	2738	7	1	2	6027	6082	
0	2739	5	1	1	6083	
0	2740	7	1	2	6028	6084	
0	2741	5	1	1	6085	
0	2742	7	1	2	6029	6086	
0	2743	5	1	1	6087	
0	2744	7	1	2	6030	6088	
0	2745	3	1	3	6355	6169	6357	
0	2746	4	1	3	6356	6170	6358	
0	2748	6	1	2	6047	2467	
0	2749	6	1	2	6043	2468	
0	2750	6	1	2	6048	2469	
0	2751	6	1	2	6044	2470	
0	2754	6	1	2	6350	2474	
0	2755	6	1	2	6348	2475	
0	2756	6	1	2	6354	2476	
0	2757	6	1	2	6352	2477	
0	2758	7	2	2	6014	2481	
0	2761	7	2	2	6050	2482	
0	2764	7	2	2	2478	1770	
0	2768	3	1	3	2486	1789	1790	
0	2769	3	1	3	2487	1797	1798	
0	2898	7	1	2	5784	2633	
0	2899	7	1	2	5788	2635	
0	2900	7	1	2	5792	2637	
0	2901	7	1	2	5796	2639	
0	2962	5	1	1	2746	
0	2966	6	1	2	2748	2749	
0	2967	6	4	2	2750	2751	
0	2973	6	5	2	2754	2755	
0	2977	6	5	2	2756	2757	
0	2980	7	1	2	6359	2143	
0	2984	5	1	1	6203	
0	2985	5	1	1	6219	
0	2986	5	1	1	6235	
0	2987	5	1	1	6251	
0	2988	5	1	1	6267	
0	2989	5	1	1	6283	
0	2990	5	1	1	6299	
0	2991	5	1	1	6315	
0	2992	5	1	1	6204	
0	2993	5	1	1	6220	
0	2994	5	1	1	6236	
0	2995	5	1	1	6252	
0	2996	5	1	1	6268	
0	2997	5	1	1	6284	
0	2998	5	1	1	6300	
0	2999	5	1	1	6316	
0	3000	5	1	1	6205	
0	3001	5	1	1	6221	
0	3002	5	1	1	6237	
0	3003	5	1	1	6253	
0	3004	5	1	1	6269	
0	3005	5	1	1	6285	
0	3006	5	1	1	6301	
0	3007	5	1	1	6317	
0	3008	5	1	1	6206	
0	3009	5	1	1	6222	
0	3010	5	1	1	6238	
0	3011	5	1	1	6254	
0	3012	5	1	1	6270	
0	3013	5	1	1	6286	
0	3014	5	1	1	6302	
0	3015	5	1	1	6318	
0	3016	5	1	1	6207	
0	3017	5	1	1	6223	
0	3018	5	1	1	6239	
0	3019	5	1	1	6255	
0	3020	5	1	1	6271	
0	3021	5	1	1	6287	
0	3022	5	1	1	6303	
0	3023	5	1	1	6319	
0	3024	5	1	1	6208	
0	3025	5	1	1	6224	
0	3026	5	1	1	6240	
0	3027	5	1	1	6256	
0	3028	5	1	1	6272	
0	3029	5	1	1	6288	
0	3030	5	1	1	6304	
0	3031	5	1	1	6320	
0	3032	5	1	1	6209	
0	3033	5	1	1	6225	
0	3034	5	1	1	6241	
0	3035	5	1	1	6257	
0	3036	5	1	1	6273	
0	3037	5	1	1	6289	
0	3038	5	1	1	6305	
0	3039	5	1	1	6321	
0	3040	5	1	1	6210	
0	3041	5	1	1	6226	
0	3042	5	1	1	6242	
0	3043	5	1	1	6258	
0	3044	5	1	1	6274	
0	3045	5	1	1	6290	
0	3046	5	1	1	6306	
0	3047	5	1	1	6322	
0	3048	5	1	1	6211	
0	3049	5	1	1	6227	
0	3050	5	1	1	6243	
0	3051	5	1	1	6259	
0	3052	5	1	1	6275	
0	3053	5	1	1	6291	
0	3054	5	1	1	6307	
0	3055	5	1	1	6323	
0	3056	5	1	1	6212	
0	3057	5	1	1	6228	
0	3058	5	1	1	6244	
0	3059	5	1	1	6260	
0	3060	5	1	1	6276	
0	3061	5	1	1	6292	
0	3062	5	1	1	6308	
0	3063	5	1	1	6324	
0	3064	5	1	1	6213	
0	3065	5	1	1	6229	
0	3066	5	1	1	6245	
0	3067	5	1	1	6261	
0	3068	5	1	1	6277	
0	3069	5	1	1	6293	
0	3070	5	1	1	6309	
0	3071	5	1	1	6325	
0	3072	5	1	1	6214	
0	3073	5	1	1	6230	
0	3074	5	1	1	6246	
0	3075	5	1	1	6262	
0	3076	5	1	1	6278	
0	3077	5	1	1	6294	
0	3078	5	1	1	6310	
0	3079	5	1	1	6326	
0	3080	5	1	1	6215	
0	3081	5	1	1	6231	
0	3082	5	1	1	6247	
0	3083	5	1	1	6263	
0	3084	5	1	1	6279	
0	3085	5	1	1	6295	
0	3086	5	1	1	6311	
0	3087	5	1	1	6327	
0	3088	5	1	1	6216	
0	3089	5	1	1	6232	
0	3090	5	1	1	6248	
0	3091	5	1	1	6264	
0	3092	5	1	1	6280	
0	3093	5	1	1	6296	
0	3094	5	1	1	6312	
0	3095	5	1	1	6328	
0	3096	5	1	1	6217	
0	3097	5	1	1	6233	
0	3098	5	1	1	6249	
0	3099	5	1	1	6265	
0	3100	5	1	1	6281	
0	3101	5	1	1	6297	
0	3102	5	1	1	6313	
0	3103	5	1	1	6329	
0	3104	5	1	1	6218	
0	3105	5	1	1	6234	
0	3106	5	1	1	6250	
0	3107	5	1	1	6266	
0	3108	5	1	1	6282	
0	3109	5	1	1	6298	
0	3110	5	1	1	6314	
0	3111	5	1	1	6330	
0	3115	5	2	1	6372	
0	3118	5	1	1	6369	
0	3119	7	2	2	2768	1674	
0	3125	5	2	1	6375	
0	3131	5	2	1	6384	
0	3134	5	1	1	6381	
0	3138	5	2	1	6393	
0	3141	5	1	1	6390	
0	3145	5	2	1	6402	
0	3148	5	1	1	6399	
0	3149	7	2	2	2769	1678	
0	3155	5	2	1	6407	
0	3161	5	2	1	6418	
0	3164	5	1	1	6415	
0	3168	5	2	1	6429	
0	3171	5	1	1	6426	
0	3172	7	4	2	6149	6366	
0	3175	7	4	2	6151	6378	
0	3178	7	4	2	6152	6387	
0	3181	7	4	2	6153	6396	
0	3184	7	4	2	6159	6412	
0	3187	7	4	2	6160	6423	
0	3190	5	1	1	6403	
0	3191	5	1	1	6408	
0	3192	5	1	1	6419	
0	3193	5	1	1	6430	
0	3194	7	1	5	6404	6409	6420	6431	1459	
3	3195	6	0	2	2745	2962	
0	3196	5	1	1	2966	
0	3206	3	1	3	2980	2145	2347	
0	3207	7	1	2	124	2984	
0	3208	7	1	2	5604	2985	
0	3209	7	1	2	5596	2986	
0	3210	7	1	2	5589	2987	
0	3211	7	1	2	5584	2988	
0	3212	7	1	2	5580	2989	
0	3213	7	1	2	5577	2990	
0	3214	7	1	2	5575	2991	
0	3215	7	1	2	5576	2992	
0	3216	7	1	2	5443	2993	
0	3217	7	1	2	5605	2994	
0	3218	7	1	2	5597	2995	
0	3219	7	1	2	5590	2996	
0	3220	7	1	2	5585	2997	
0	3221	7	1	2	5581	2998	
0	3222	7	1	2	5578	2999	
0	3223	7	1	2	5579	3000	
0	3224	7	1	2	5462	3001	
0	3225	7	1	2	5444	3002	
0	3226	7	1	2	5606	3003	
0	3227	7	1	2	5598	3004	
0	3228	7	1	2	5591	3005	
0	3229	7	1	2	5586	3006	
0	3230	7	1	2	5582	3007	
0	3231	7	1	2	5583	3008	
0	3232	7	1	2	5482	3009	
0	3233	7	1	2	5463	3010	
0	3234	7	1	2	5445	3011	
0	3235	7	1	2	5607	3012	
0	3236	7	1	2	5599	3013	
0	3237	7	1	2	5592	3014	
0	3238	7	1	2	5587	3015	
0	3239	7	1	2	5588	3016	
0	3240	7	1	2	5499	3017	
0	3241	7	1	2	5483	3018	
0	3242	7	1	2	5464	3019	
0	3243	7	1	2	5446	3020	
0	3244	7	1	2	5608	3021	
0	3245	7	1	2	5600	3022	
0	3246	7	1	2	5593	3023	
0	3247	7	1	2	5594	3024	
0	3248	7	1	2	5516	3025	
0	3249	7	1	2	5500	3026	
0	3250	7	1	2	5484	3027	
0	3251	7	1	2	5465	3028	
0	3252	7	1	2	5447	3029	
0	3253	7	1	2	5609	3030	
0	3254	7	1	2	5601	3031	
0	3255	7	1	2	5602	3032	
0	3256	7	1	2	5535	3033	
0	3257	7	1	2	5517	3034	
0	3258	7	1	2	5501	3035	
0	3259	7	1	2	5485	3036	
0	3260	7	1	2	5466	3037	
0	3261	7	1	2	5448	3038	
0	3262	7	1	2	5610	3039	
0	3263	7	1	2	5611	3040	
0	3264	7	1	2	5553	3041	
0	3265	7	1	2	5536	3042	
0	3266	7	1	2	5518	3043	
0	3267	7	1	2	5502	3044	
0	3268	7	1	2	5486	3045	
0	3269	7	1	2	5467	3046	
0	3270	7	1	2	5449	3047	
0	3271	7	1	2	5722	3048	
0	3272	7	1	2	5468	3049	
0	3273	7	1	2	5487	3050	
0	3274	7	1	2	5503	3051	
0	3275	7	1	2	5519	3052	
0	3276	7	1	2	5537	3053	
0	3277	7	1	2	5554	3054	
0	3278	7	1	2	5568	3055	
0	3279	7	1	2	5731	3056	
0	3280	7	1	2	5488	3057	
0	3281	7	1	2	5504	3058	
0	3282	7	1	2	5520	3059	
0	3283	7	1	2	5538	3060	
0	3284	7	1	2	5555	3061	
0	3285	7	1	2	5569	3062	
0	3286	7	1	2	5723	3063	
0	3287	7	1	2	5739	3064	
0	3288	7	1	2	5505	3065	
0	3289	7	1	2	5521	3066	
0	3290	7	1	2	5539	3067	
0	3291	7	1	2	5556	3068	
0	3292	7	1	2	5570	3069	
0	3293	7	1	2	5724	3070	
0	3294	7	1	2	5732	3071	
0	3295	7	1	2	5745	3072	
0	3296	7	1	2	5522	3073	
0	3297	7	1	2	5540	3074	
0	3298	7	1	2	5557	3075	
0	3299	7	1	2	5571	3076	
0	3300	7	1	2	5725	3077	
0	3301	7	1	2	5733	3078	
0	3302	7	1	2	5740	3079	
0	3303	7	1	2	5750	3080	
0	3304	7	1	2	5541	3081	
0	3305	7	1	2	5558	3082	
0	3306	7	1	2	5572	3083	
0	3307	7	1	2	5726	3084	
0	3308	7	1	2	5734	3085	
0	3309	7	1	2	5741	3086	
0	3310	7	1	2	5746	3087	
0	3311	7	1	2	5754	3088	
0	3312	7	1	2	5559	3089	
0	3313	7	1	2	5573	3090	
0	3314	7	1	2	5727	3091	
0	3315	7	1	2	5735	3092	
0	3316	7	1	2	5742	3093	
0	3317	7	1	2	5747	3094	
0	3318	7	1	2	5751	3095	
0	3319	7	1	2	5757	3096	
0	3320	7	1	2	5574	3097	
0	3321	7	1	2	5728	3098	
0	3322	7	1	2	5736	3099	
0	3323	7	1	2	5743	3100	
0	3324	7	1	2	5748	3101	
0	3325	7	1	2	5752	3102	
0	3326	7	1	2	5755	3103	
0	3327	7	1	2	329	3104	
0	3328	7	1	2	5729	3105	
0	3329	7	1	2	5737	3106	
0	3330	7	1	2	5744	3107	
0	3331	7	1	2	5749	3108	
0	3332	7	1	2	5753	3109	
0	3333	7	1	2	5756	3110	
0	3334	7	1	2	5758	3111	
0	3383	7	1	5	3190	3191	3192	3193	5623	
0	3387	7	1	2	3196	1736	
0	3388	7	1	2	6449	2149	
0	3389	7	1	2	6444	1737	
0	3390	4	1	8	3207	3208	3209	3210	3211	3212	3213	3214	
0	3391	4	1	8	3215	3216	3217	3218	3219	3220	3221	3222	
0	3392	4	1	8	3223	3224	3225	3226	3227	3228	3229	3230	
0	3393	4	1	8	3231	3232	3233	3234	3235	3236	3237	3238	
0	3394	4	1	8	3239	3240	3241	3242	3243	3244	3245	3246	
0	3395	4	1	8	3247	3248	3249	3250	3251	3252	3253	3254	
0	3396	4	1	8	3255	3256	3257	3258	3259	3260	3261	3262	
0	3397	4	1	8	3263	3264	3265	3266	3267	3268	3269	3270	
0	3398	4	1	8	3271	3272	3273	3274	3275	3276	3277	3278	
0	3399	4	1	8	3279	3280	3281	3282	3283	3284	3285	3286	
0	3400	4	1	8	3287	3288	3289	3290	3291	3292	3293	3294	
0	3401	4	1	8	3295	3296	3297	3298	3299	3300	3301	3302	
0	3402	4	1	8	3303	3304	3305	3306	3307	3308	3309	3310	
0	3403	4	1	8	3311	3312	3313	3314	3315	3316	3317	3318	
0	3404	4	1	8	3319	3320	3321	3322	3323	3324	3325	3326	
0	3405	4	1	8	3327	3328	3329	3330	3331	3332	3333	3334	
0	3406	7	1	2	3206	2641	
0	3407	7	2	3	5613	6367	6373	
0	3410	7	2	3	5624	6368	6454	
0	3413	7	1	3	5634	6370	6455	
0	3414	7	1	3	5646	6371	6374	
0	3415	3	3	3	6456	6135	6189	
0	3419	4	3	3	6457	6136	6190	
0	3423	7	2	3	5614	6379	6385	
0	3426	7	2	3	5625	6380	6460	
0	3429	7	1	3	5635	6382	6461	
0	3430	7	1	3	5647	6383	6386	
0	3431	7	2	3	5615	6388	6394	
0	3434	7	2	3	5626	6389	6462	
0	3437	7	1	3	5636	6391	6463	
0	3438	7	1	3	5648	6392	6395	
0	3439	7	2	3	5616	6397	6405	
0	3442	7	2	3	5627	6398	6464	
0	3445	7	1	3	5637	6400	6465	
0	3446	7	1	3	5649	6401	6406	
0	3447	3	3	3	6466	6143	6197	
0	3451	4	3	3	6467	6144	6198	
0	3455	7	2	3	5617	6413	6421	
0	3458	7	2	3	5628	6414	6470	
0	3461	7	1	3	5638	6416	6471	
0	3462	7	1	3	5650	6417	6422	
0	3463	7	2	3	5618	6424	6432	
0	3466	7	2	3	5629	6425	6472	
0	3469	7	1	3	5639	6427	6473	
0	3470	7	1	3	5651	6428	6433	
0	3471	3	1	2	3194	3383	
0	3534	4	1	2	3387	2350	
0	3535	3	1	3	3388	2151	2351	
0	3536	4	1	2	3389	1966	
0	3537	7	1	2	3390	2209	
0	3538	7	1	2	3398	2210	
0	3539	7	1	2	3391	1842	
0	3540	7	1	2	3399	5419	
0	3541	7	1	2	3392	1843	
0	3542	7	1	2	3400	5420	
0	3543	7	1	2	3393	1844	
0	3544	7	1	2	3401	5421	
0	3545	7	1	2	3394	1845	
0	3546	7	1	2	3402	5422	
0	3547	7	1	2	3395	1846	
0	3548	7	1	2	3403	5423	
0	3549	7	1	2	3396	1847	
0	3550	7	1	2	3404	5424	
0	3551	7	1	2	3397	1848	
0	3552	7	1	2	3405	5425	
0	3557	3	1	3	3413	3414	3118	
0	3568	3	1	3	3429	3430	3134	
0	3573	3	1	3	3437	3438	3141	
0	3578	3	1	3	3445	3446	3148	
0	3589	3	1	3	3461	3462	3164	
0	3594	3	1	3	3469	3470	3171	
0	3605	7	1	2	3471	2728	
0	3626	5	1	1	6440	
0	3627	5	1	1	6360	
0	3628	5	1	1	6445	
0	3629	5	1	1	6446	
0	3630	5	1	1	6441	
0	3631	5	1	1	6361	
0	3632	7	1	2	3536	2152	
0	3633	7	1	2	3534	2155	
0	3634	3	1	3	3537	3538	2398	
0	3635	3	1	2	3539	3540	
0	3636	3	1	2	3541	3542	
0	3637	3	1	2	3543	3544	
0	3638	3	1	2	3545	3546	
0	3639	3	1	2	3547	3548	
0	3640	3	1	2	3549	3550	
0	3641	3	1	2	3551	3552	
0	3642	7	1	2	3535	2643	
0	3643	3	1	2	6498	6500	
0	3644	4	1	2	6499	6501	
0	3645	7	2	3	5619	6502	6376	
0	3648	7	2	3	5630	6503	6458	
0	3651	7	1	3	5640	6505	6459	
0	3652	7	1	3	5652	6506	6377	
0	3653	5	1	1	6507	
0	3654	3	2	2	6508	6510	
0	3657	4	1	2	6509	6511	
0	3658	3	2	2	6512	6514	
0	3661	4	1	2	6513	6515	
0	3662	3	1	2	6516	6518	
0	3663	4	1	2	6517	6519	
0	3664	7	2	3	5620	6520	6410	
0	3667	7	2	3	5631	6521	6468	
0	3670	7	1	3	5641	6523	6469	
0	3671	7	1	3	5653	6524	6411	
0	3672	5	1	1	6525	
0	3673	3	2	2	6526	6528	
0	3676	4	1	2	6527	6529	
0	3677	3	2	2	6530	6532	
0	3680	4	1	2	6531	6533	
0	3681	5	1	1	6474	
0	3682	7	4	2	6150	6504	
0	3685	5	1	1	6478	
0	3686	5	1	1	6479	
0	3687	5	1	1	6482	
0	3688	5	1	1	6483	
0	3689	5	1	1	6486	
0	3690	7	4	2	6161	6522	
0	3693	5	1	1	6490	
0	3694	5	1	1	6494	
0	3695	5	1	1	6495	
0	3696	5	1	1	6491	
0	3703	5	1	1	6475	
0	3704	5	1	1	6487	
0	3705	6	1	2	6362	3630	
0	3706	6	1	2	6442	3631	
0	3707	6	1	2	6363	3626	
0	3708	6	1	2	6443	3627	
0	3711	3	1	3	3632	2352	2353	
0	3712	3	1	3	3633	2354	2355	
0	3713	7	1	2	3634	2632	
0	3714	7	1	2	3635	2634	
0	3715	7	1	2	3636	2636	
0	3716	7	1	2	3637	2638	
0	3717	7	1	2	3638	2640	
0	3718	7	1	2	3639	2642	
0	3719	7	1	2	3640	2644	
0	3720	7	1	2	3641	2646	
0	3721	7	8	2	3644	3557	
0	3731	3	1	3	3651	3652	3653	
0	3734	7	6	2	3657	3568	
0	3740	7	5	2	3661	3573	
0	3743	7	8	2	3663	3578	
0	3753	3	1	3	3670	3671	3672	
0	3756	7	6	2	3676	3589	
0	3762	7	5	2	3680	3594	
0	3765	5	1	1	3643	
0	3766	5	1	1	3662	
0	3773	6	1	2	3705	3706	
0	3774	6	1	2	3707	3708	
0	3775	6	1	2	6450	3628	
0	3776	5	1	1	6451	
0	3777	6	1	2	6452	3629	
0	3778	5	1	1	6453	
0	3779	7	1	2	3712	2645	
0	3780	7	1	2	3711	2647	
0	3786	3	2	2	6534	6536	
0	3789	4	1	2	6535	6537	
0	3800	3	2	2	6542	6544	
0	3803	4	1	2	6543	6545	
0	3809	7	2	2	6538	6155	
0	3812	7	3	2	6540	6156	
0	3815	7	2	2	6546	6162	
0	3818	7	4	2	6548	6163	
3	3833	6	0	2	3773	3774	
0	3834	6	1	2	6447	3776	
0	3835	6	1	2	6448	3778	
0	3838	7	7	2	3789	3731	
0	3845	7	7	2	3803	3753	
0	3884	6	1	2	3775	3834	
0	3885	6	1	2	3777	3835	
0	3894	6	1	2	6558	6596	
0	3895	6	1	2	6577	6598	
0	3898	5	1	1	6550	
0	3899	5	1	1	6551	
0	3906	5	1	1	6554	
0	3911	5	1	1	6555	
0	3912	7	1	2	6597	1912	
0	3916	7	1	2	6599	6157	
0	3920	5	1	1	6600	
0	3924	5	1	1	3884	
0	3925	5	1	1	3885	
0	3926	7	4	4	6559	6611	6566	6572	
0	3930	6	1	3	6560	6612	6539	
0	3931	6	1	4	6541	6613	6567	6561	
0	3932	7	2	4	6578	6618	6585	6591	
0	3935	6	1	3	6579	6619	6547	
0	3936	6	1	4	6549	6620	6586	6580	
0	3947	5	1	1	3912	
0	3948	5	1	1	3916	
3	3987	6	0	2	3924	3925	
0	3992	6	2	4	3765	3894	3930	3931	
0	3996	6	2	4	3766	3895	3935	3936	
0	4013	5	1	1	6607	
3	4028	7	0	2	6629	6625	
0	4029	6	1	2	6562	3681	
0	4030	6	1	2	6568	3686	
0	4031	6	1	2	6573	3688	
0	4032	6	1	2	6581	3689	
0	4033	6	1	2	6587	3693	
0	4034	6	1	2	6592	3695	
0	4042	5	1	1	6563	
0	4043	5	1	1	6569	
0	4044	6	1	2	6570	3685	
0	4045	5	1	1	6571	
0	4046	5	1	1	6574	
0	4047	6	1	2	6575	3687	
0	4048	5	1	1	6576	
0	4049	5	1	1	6582	
0	4050	5	1	1	6588	
0	4051	5	1	1	6593	
0	4052	6	1	2	6594	3694	
0	4053	5	1	1	6595	
0	4054	5	1	1	6589	
0	4055	6	1	2	6590	3696	
0	4056	7	1	2	6630	6158	
0	4057	5	1	1	6564	
0	4058	6	1	2	6565	3703	
0	4065	5	1	1	6583	
0	4066	6	1	2	6584	3704	
0	4073	6	1	2	6626	6633	
0	4074	5	1	1	6631	
0	4075	6	1	2	6476	4042	
0	4076	6	1	2	6480	4045	
0	4077	6	1	2	6484	4048	
0	4078	6	1	2	6488	4049	
0	4079	6	1	2	6492	4050	
0	4080	6	1	2	6496	4053	
0	4085	6	1	2	6481	4043	
0	4086	6	1	2	6485	4046	
0	4088	6	1	2	6497	4051	
0	4090	6	1	2	6493	4054	
0	4091	7	9	2	6634	6164	
0	4094	3	6	2	3605	4056	
0	4098	6	1	2	6477	4057	
0	4101	6	1	2	6489	4065	
0	4104	7	1	2	4073	4074	
0	4105	6	1	2	4075	4029	
0	4106	6	1	2	6614	3899	
0	4107	6	1	2	4076	4030	
0	4108	6	1	2	4077	4031	
0	4109	6	1	2	4078	4032	
0	4110	6	1	2	6621	3906	
0	4111	6	1	2	4079	4033	
0	4112	6	1	2	4080	4034	
0	4113	5	1	1	6615	
0	4114	6	1	2	6616	3898	
0	4115	5	1	1	6617	
0	4116	6	8	2	4085	4044	
0	4119	6	8	2	4086	4047	
0	4122	5	1	1	6622	
0	4123	6	5	2	4088	4052	
0	4126	5	1	1	6623	
0	4127	6	1	2	6624	3911	
0	4128	6	6	2	4090	4055	
0	4139	6	2	2	4098	4058	
0	4142	6	2	2	4101	4066	
3	4145	5	0	1	4104	
0	4146	5	1	1	4105	
0	4147	6	1	2	6552	4115	
0	4148	5	1	1	4107	
0	4149	5	1	1	4108	
0	4150	5	1	1	4109	
0	4151	6	1	2	6556	4122	
0	4152	5	1	1	4111	
0	4153	5	1	1	4112	
0	4154	6	1	2	6553	4113	
0	4161	6	1	2	6557	4126	
0	4186	7	2	2	5760	6644	
0	4189	7	1	2	4146	2230	
0	4190	6	1	2	4147	4106	
0	4191	7	1	2	4148	2232	
0	4192	7	1	2	4149	2233	
0	4193	7	1	2	4150	2234	
0	4194	6	1	2	4151	4110	
0	4195	7	1	2	4152	2236	
0	4196	7	1	2	4153	2237	
0	4197	6	6	2	4154	4114	
0	4218	6	5	2	4161	4127	
0	4238	7	1	2	6671	6608	
0	4239	5	1	1	6677	
0	4241	5	1	1	6679	
0	4242	7	4	2	5761	6666	
0	4251	4	1	3	3713	4189	2898	
0	4252	5	1	1	4190	
0	4253	4	1	3	3715	4191	2900	
0	4254	4	1	3	3716	4192	2901	
0	4255	4	1	3	3717	4193	3406	
0	4256	5	1	1	4194	
0	4257	4	1	3	3719	4195	3779	
0	4258	4	1	3	3720	4196	3780	
0	4283	7	1	2	6635	6627	
0	4284	7	3	2	6645	6628	
0	4287	3	5	2	6605	4238	
0	4291	5	1	1	6681	
0	4295	5	1	1	6636	
0	4299	5	1	1	6637	
0	4303	7	1	2	4252	2231	
0	4304	7	1	2	4256	2235	
0	4310	3	5	2	6632	4283	
0	4316	7	1	3	6646	6658	6650	
0	4317	7	1	2	6647	6659	
0	4318	7	1	3	6667	6672	6689	
0	4319	7	2	2	6668	6673	
0	4322	7	1	2	6638	6660	
0	4325	6	1	2	6651	6602	
0	4326	6	1	3	6652	6661	6639	
0	4327	6	1	2	6690	6606	
0	4328	6	1	3	6691	6674	6609	
0	4329	6	1	2	6675	4013	
0	4330	5	1	1	6676	
0	4331	7	2	3	5762	6648	4295	
0	4335	7	2	2	4251	2730	
0	4338	7	2	2	4253	2734	
0	4341	7	2	2	4254	2736	
0	4344	7	2	2	4255	2738	
0	4347	7	2	2	4257	2742	
0	4350	7	2	2	4258	2744	
0	4371	7	2	2	6669	6670	
0	4376	4	1	3	3714	4303	2899	
0	4377	4	1	3	3718	4304	3642	
0	4387	7	4	2	5763	4317	
0	4390	7	4	2	5764	4318	
0	4393	6	1	2	6610	4330	
0	4416	6	2	3	3920	4325	4326	
0	4421	3	2	2	6603	4322	
0	4427	6	2	3	3948	4327	4328	
0	4435	7	2	2	5765	4316	
0	4442	3	1	2	6713	6640	
0	4443	7	3	4	6649	6683	6653	6662	
0	4446	6	1	2	6684	6601	
0	4447	6	1	3	6685	6654	6604	
0	4448	6	1	4	6686	6655	6663	6641	
0	4452	5	1	1	6656	
0	4458	6	4	2	4329	4393	
0	4461	5	1	1	6694	
0	4462	5	1	1	6695	
0	4463	6	1	2	6727	1460	
0	4464	5	1	1	6728	
0	4468	4	5	2	6714	6642	
0	4472	7	2	2	4376	2732	
0	4475	7	2	2	4377	2740	
0	4484	5	1	1	6687	
0	4486	5	1	1	6664	
0	4487	6	1	2	6665	4299	
0	4491	5	1	1	6692	
0	4493	7	2	2	5766	6711	
0	4496	5	1	1	6701	
0	4497	7	1	2	6702	6703	
0	4498	7	2	2	4442	1769	
0	4503	6	4	4	3947	4446	4447	4448	
0	4506	5	1	1	6698	
0	4507	5	1	1	6743	
0	4508	5	1	1	6739	
0	4509	6	1	2	6740	4452	
0	4510	5	1	1	6741	
0	4511	6	1	2	6742	4241	
0	4515	6	1	2	5767	4464	
0	4526	5	1	1	6737	
0	4527	6	1	2	6738	4484	
0	4528	6	1	2	6643	4486	
0	4529	5	1	1	6704	
0	4530	6	1	2	6705	4491	
0	4545	7	1	3	5768	6712	4496	
0	4549	7	4	2	5769	6745	
0	4552	6	1	2	6657	4508	
0	4555	6	1	2	6680	4510	
0	4558	5	1	1	6761	
0	4559	6	2	2	4463	4515	
0	4562	5	1	1	6706	
0	4563	7	1	2	6707	6708	
0	4568	5	1	1	6709	
0	4572	6	1	2	6688	4526	
0	4573	6	1	2	6693	4529	
0	4576	6	2	2	4487	4528	
0	4587	3	1	3	6434	6763	6436	
0	4588	4	1	3	6435	6764	6437	
3	4589	3	0	2	4545	4497	
0	4593	6	4	2	4552	4509	
0	4596	5	1	1	6729	
0	4597	5	1	1	6730	
0	4599	6	4	2	4555	4511	
0	4602	5	1	1	6733	
0	4603	5	1	1	6734	
0	4608	7	1	3	5770	6699	4562	
0	4619	6	2	2	4572	4527	
0	4623	6	2	2	4573	4530	
0	4628	5	1	1	4588	
0	4629	6	1	2	6746	4506	
0	4630	5	1	1	6747	
0	4635	5	1	1	6775	
0	4636	6	1	2	6776	4291	
0	4640	5	1	1	6748	
0	4641	6	1	2	6749	4461	
0	4642	5	1	1	6750	
0	4643	6	1	2	6751	4462	
0	4644	4	5	2	4608	4563	
0	4647	7	2	2	6773	2128	
0	4650	7	2	2	6774	2743	
3	4667	7	0	2	4587	4628	
0	4668	6	1	2	6700	4630	
0	4669	5	1	1	6765	
0	4670	6	1	2	6766	4239	
0	4673	5	1	1	6785	
0	4674	6	1	2	6786	4507	
0	4675	6	1	2	6682	4635	
0	4676	5	1	1	6787	
0	4677	6	1	2	6788	4558	
0	4678	6	1	2	6696	4640	
0	4679	6	1	2	6697	4642	
0	4687	5	1	1	6767	
0	4688	6	1	2	6768	4568	
0	4704	6	1	2	4629	4668	
0	4705	6	1	2	6678	4669	
0	4706	5	1	1	6769	
0	4707	5	1	1	6770	
0	4708	6	1	2	6744	4673	
0	4711	6	2	2	4675	4636	
0	4716	6	1	2	6762	4676	
0	4717	6	3	2	4678	4641	
0	4721	6	1	2	4679	4643	
0	4726	5	1	1	6752	
0	4727	3	3	3	6794	6796	6725	
0	4730	4	2	3	6795	6797	6726	
0	4733	6	1	2	6710	4687	
0	4740	6	4	2	4705	4670	
0	4743	6	4	2	4708	4674	
0	4747	5	1	1	6777	
0	4748	6	1	2	6778	4596	
0	4749	5	1	1	6779	
0	4750	6	1	2	6780	4597	
0	4753	5	1	1	6781	
0	4754	6	1	2	6782	4602	
0	4755	5	1	1	6783	
0	4756	6	1	2	6784	4603	
0	4757	6	4	2	4716	4677	
0	4769	6	2	2	4733	4688	
0	4772	7	2	2	5771	4704	
0	4775	5	2	1	4721	
0	4778	5	1	1	6806	
0	4786	6	1	2	6731	4747	
0	4787	6	1	2	6732	4749	
0	4788	6	1	2	6735	4753	
0	4789	6	1	2	6736	4755	
0	4794	7	2	2	6798	2124	
0	4797	7	2	2	6799	2735	
0	4800	7	2	2	6800	2127	
0	4808	7	2	2	6801	6753	
3	4815	7	0	2	6803	4778	
0	4816	5	1	1	6820	
0	4817	5	1	1	6822	
0	4818	6	3	2	4786	4748	
0	4822	6	1	2	4787	4750	
0	4823	6	2	2	4788	4754	
0	4826	6	1	2	4789	4756	
0	4829	6	1	2	6824	4726	
0	4830	5	1	1	6825	
0	4831	7	2	2	6812	2122	
0	4838	7	2	2	6816	2126	
0	4859	6	1	2	6823	4816	
0	4860	6	1	2	6821	4817	
0	4868	5	1	1	4826	
0	4870	5	1	1	6789	
0	4872	5	1	1	6832	
0	4873	6	1	2	6754	4830	
0	4876	3	5	3	6826	6828	6719	
0	4880	4	2	3	6827	6829	6720	
0	4885	5	1	1	6804	
0	4889	5	2	1	4822	
0	4895	6	1	2	4859	4860	
0	4896	5	1	1	6808	
0	4897	6	1	2	6809	4706	
0	4898	5	1	1	6810	
0	4899	6	1	2	6811	4707	
0	4900	4	1	2	4868	6755	
0	4901	7	1	4	6802	6817	6837	6756	
0	4902	5	1	1	6813	
0	4904	5	1	1	6818	
0	4905	6	1	2	6819	4872	
0	4906	6	1	2	4873	4829	
0	4907	7	2	2	6834	2123	
0	4913	7	2	2	6838	2125	
0	4916	7	2	2	6835	6790	
0	4920	5	1	1	6848	
0	4921	7	2	2	4895	2184	
0	4924	6	1	2	6771	4896	
0	4925	6	1	2	6772	4898	
0	4926	3	1	2	4900	4901	
0	4928	6	1	2	6850	4870	
0	4929	5	1	1	6851	
0	4930	6	1	2	6833	4904	
0	4931	5	1	1	4906	
3	4944	7	0	2	6843	4920	
0	4946	6	2	2	4924	4897	
0	4949	6	1	2	4925	4899	
0	4950	6	1	2	6856	4902	
0	4951	5	1	1	6857	
0	4952	6	1	2	6791	4929	
0	4953	6	1	2	4930	4905	
0	4954	7	2	2	4926	2737	
0	4957	7	2	2	4931	2741	
0	4964	3	1	3	6438	6364	6858	
0	4965	4	1	3	6439	6365	6859	
0	4968	5	1	1	4949	
0	4969	6	1	2	6814	4951	
0	4970	6	1	2	4952	4928	
0	4973	7	2	2	4953	2739	
0	4978	5	1	1	6844	
0	4979	5	1	1	6845	
0	4980	5	1	1	4965	
0	4981	4	1	2	4968	6792	
0	4982	7	1	4	6836	6815	6860	6793	
0	4983	6	1	2	4950	4969	
0	4984	5	1	1	4970	
0	4985	7	2	2	6861	2121	
0	4988	3	3	3	6854	6862	6721	
0	4991	4	2	3	6855	6863	6722	
0	4996	3	3	3	6830	6864	6723	
0	4999	4	2	3	6831	6865	6724	
3	5002	7	0	2	4964	4980	
0	5007	3	1	2	4981	4982	
0	5010	7	2	2	4983	2731	
0	5013	7	2	2	4984	2733	
0	5018	3	3	3	6841	6866	6759	
0	5021	4	2	3	6842	6867	6760	
0	5026	5	1	1	6873	
0	5029	5	1	1	6878	
0	5030	7	2	2	5007	2729	
3	5045	7	0	2	6870	5026	
0	5046	5	1	1	6887	
3	5047	7	0	2	6875	5029	
0	5050	3	5	3	6839	6880	6757	
0	5055	4	2	3	6840	6881	6758	
0	5058	3	5	3	6852	6882	6717	
0	5061	4	2	3	6853	6883	6718	
0	5066	7	2	4	6807	6879	6888	6874	
3	5078	7	0	2	6884	5046	
0	5080	3	5	3	6868	6889	6715	
0	5085	4	2	3	6869	6890	6716	
0	5094	6	1	2	6876	4885	
0	5095	5	1	1	6877	
0	5097	5	1	1	6871	
3	5102	7	0	2	6891	6892	
0	5103	5	1	1	6903	
0	5108	6	1	2	6805	5095	
0	5109	5	1	1	6885	
0	5110	6	1	2	6886	5097	
0	5114	7	4	2	6893	6007	
3	5120	7	0	2	6907	6908	
3	5121	7	0	2	6898	5103	
0	5122	6	4	2	5094	5108	
0	5125	6	1	2	6872	5109	
0	5128	7	4	2	6008	6909	
0	5133	7	2	4	6849	6904	6896	6912	
0	5136	7	1	3	6897	6913	6011	
0	5145	6	4	2	5125	5110	
0	5159	5	1	1	6894	
0	5166	7	1	2	6905	6926	
0	5173	7	1	2	6906	6927	
0	5182	5	1	1	6910	
0	5183	6	1	2	6911	5159	
3	5192	5	0	1	5166	
0	5193	4	1	2	5136	5173	
0	5196	6	1	2	6899	4978	
0	5197	5	1	1	6900	
0	5198	6	1	2	6901	4979	
0	5199	5	1	1	6902	
0	5201	5	1	1	6914	
0	5203	5	1	1	6915	
0	5212	6	1	2	6895	5182	
0	5215	7	1	2	5661	5193	
0	5217	5	1	1	6918	
0	5219	5	1	1	6919	
0	5220	6	1	2	6846	5197	
0	5221	6	1	2	6847	5199	
0	5222	5	1	1	6922	
0	5223	6	1	2	6923	5201	
0	5224	6	1	2	6924	5203	
0	5225	5	1	1	6925	
0	5228	6	2	2	5183	5212	
3	5231	5	0	1	5215	
0	5232	6	1	2	6928	5217	
0	5233	5	1	1	6929	
0	5234	6	1	2	6930	5219	
0	5235	5	1	1	6931	
0	5236	6	4	2	5196	5220	
0	5240	6	1	2	5198	5221	
0	5242	6	1	2	6916	5222	
0	5243	6	1	2	6917	5225	
0	5245	6	1	2	6920	5233	
0	5246	6	1	2	6921	5235	
0	5250	5	2	1	5240	
0	5253	5	1	1	6932	
0	5254	6	2	2	5242	5223	
0	5257	6	1	2	5243	5224	
0	5258	6	4	2	5232	5245	
0	5261	6	1	2	5234	5246	
0	5266	5	2	1	5257	
0	5277	7	1	3	6934	6940	6343	
0	5278	7	1	3	6938	6941	6345	
0	5279	5	4	1	5261	
0	5283	5	1	1	6935	
0	5284	6	1	2	6936	5253	
0	5285	7	1	3	6937	6946	6346	
0	5286	7	1	3	6939	6947	6344	
0	5295	6	1	2	6933	5283	
0	5298	3	4	4	5277	5285	5278	5286	
0	5309	6	4	2	5295	5284	
0	5312	5	1	1	6942	
0	5313	5	1	1	6943	
0	5322	5	1	1	6948	
0	5323	5	1	1	6949	
0	5340	6	1	2	6952	5323	
0	5341	6	1	2	6953	5322	
0	5344	5	1	1	6954	
0	5345	5	1	1	6955	
0	5348	6	1	2	6956	5313	
0	5349	6	1	2	6957	5312	
0	5350	6	1	2	6950	5345	
0	5351	6	1	2	6951	5344	
0	5352	5	1	1	6958	
0	5353	5	1	1	6959	
0	5354	6	1	2	6944	5353	
0	5355	6	1	2	6945	5352	
0	5356	6	1	2	5350	5340	
0	5357	6	1	2	5351	5341	
0	5358	6	1	2	5348	5354	
0	5359	6	1	2	5349	5355	
3	5360	7	0	2	5356	5357	
3	5361	6	0	2	5358	5359	
2	5362	1	1			
2	5363	1	1			
2	5364	1	1			
2	5365	1	1			
2	5366	1	1			
2	5367	1	1			
2	5368	1	1			
2	5369	1	1			
2	5370	1	1			
2	5371	1	1			
2	5372	1	1			
2	5373	1	1			
2	5374	1	1			
2	5375	1	1			
2	5376	1	1			
2	5377	1	1			
2	5378	1	1			
2	5379	1	1			
2	5380	1	13			
2	5381	1	13			
2	5382	1	13			
2	5383	1	13			
2	5384	1	13			
2	5385	1	13			
2	5386	1	13			
2	5387	1	13			
2	5388	1	13			
2	5389	1	20			
2	5390	1	20			
2	5391	1	20			
2	5392	1	20			
2	5393	1	20			
2	5394	1	20			
2	5395	1	20			
2	5396	1	20			
2	5397	1	20			
2	5398	1	20			
2	5399	1	20			
2	5400	1	20			
2	5401	1	20			
2	5402	1	20			
2	5403	1	20			
2	5404	1	33			
2	5405	1	33			
2	5406	1	33			
2	5407	1	33			
2	5408	1	33			
2	5409	1	33			
2	5410	1	33			
2	5411	1	33			
2	5412	1	33			
2	5413	1	33			
2	5414	1	33			
2	5415	1	33			
2	5416	1	33			
2	5417	1	33			
2	5418	1	33			
2	5419	1	33			
2	5420	1	33			
2	5421	1	33			
2	5422	1	33			
2	5423	1	33			
2	5424	1	33			
2	5425	1	33			
2	5426	1	41			
2	5427	1	41			
2	5428	1	41			
2	5429	1	45			
2	5430	1	45			
2	5431	1	45			
2	5432	1	45			
2	5433	1	45			
2	5434	1	50			
2	5435	1	50			
2	5436	1	50			
2	5437	1	50			
2	5438	1	50			
2	5439	1	50			
2	5440	1	50			
2	5441	1	50			
2	5442	1	50			
2	5443	1	50			
2	5444	1	50			
2	5445	1	50			
2	5446	1	50			
2	5447	1	50			
2	5448	1	50			
2	5449	1	50			
2	5450	1	58			
2	5451	1	58			
2	5452	1	58			
2	5453	1	58			
2	5454	1	58			
2	5455	1	58			
2	5456	1	58			
2	5457	1	58			
2	5458	1	58			
2	5459	1	58			
2	5460	1	58			
2	5461	1	58			
2	5462	1	58			
2	5463	1	58			
2	5464	1	58			
2	5465	1	58			
2	5466	1	58			
2	5467	1	58			
2	5468	1	58			
2	5469	1	68			
2	5470	1	68			
2	5471	1	68			
2	5472	1	68			
2	5473	1	68			
2	5474	1	68			
2	5475	1	68			
2	5476	1	68			
2	5477	1	68			
2	5478	1	68			
2	5479	1	68			
2	5480	1	68			
2	5481	1	68			
2	5482	1	68			
2	5483	1	68			
2	5484	1	68			
2	5485	1	68			
2	5486	1	68			
2	5487	1	68			
2	5488	1	68			
2	5489	1	77			
2	5490	1	77			
2	5491	1	77			
2	5492	1	77			
2	5493	1	77			
2	5494	1	77			
2	5495	1	77			
2	5496	1	77			
2	5497	1	77			
2	5498	1	77			
2	5499	1	77			
2	5500	1	77			
2	5501	1	77			
2	5502	1	77			
2	5503	1	77			
2	5504	1	77			
2	5505	1	77			
2	5506	1	87			
2	5507	1	87			
2	5508	1	87			
2	5509	1	87			
2	5510	1	87			
2	5511	1	87			
2	5512	1	87			
2	5513	1	87			
2	5514	1	87			
2	5515	1	87			
2	5516	1	87			
2	5517	1	87			
2	5518	1	87			
2	5519	1	87			
2	5520	1	87			
2	5521	1	87			
2	5522	1	87			
2	5523	1	97			
2	5524	1	97			
2	5525	1	97			
2	5526	1	97			
2	5527	1	97			
2	5528	1	97			
2	5529	1	97			
2	5530	1	97			
2	5531	1	97			
2	5532	1	97			
2	5533	1	97			
2	5534	1	97			
2	5535	1	97			
2	5536	1	97			
2	5537	1	97			
2	5538	1	97			
2	5539	1	97			
2	5540	1	97			
2	5541	1	97			
2	5542	1	107			
2	5543	1	107			
2	5544	1	107			
2	5545	1	107			
2	5546	1	107			
2	5547	1	107			
2	5548	1	107			
2	5549	1	107			
2	5550	1	107			
2	5551	1	107			
2	5552	1	107			
2	5553	1	107			
2	5554	1	107			
2	5555	1	107			
2	5556	1	107			
2	5557	1	107			
2	5558	1	107			
2	5559	1	107			
2	5560	1	116			
2	5561	1	116			
2	5562	1	116			
2	5563	1	116			
2	5564	1	116			
2	5565	1	116			
2	5566	1	116			
2	5567	1	116			
2	5568	1	116			
2	5569	1	116			
2	5570	1	116			
2	5571	1	116			
2	5572	1	116			
2	5573	1	116			
2	5574	1	116			
2	5575	1	125			
2	5576	1	125			
2	5577	1	128			
2	5578	1	128			
2	5579	1	128			
2	5580	1	132			
2	5581	1	132			
2	5582	1	132			
2	5583	1	132			
2	5584	1	137			
2	5585	1	137			
2	5586	1	137			
2	5587	1	137			
2	5588	1	137			
2	5589	1	143			
2	5590	1	143			
2	5591	1	143			
2	5592	1	143			
2	5593	1	143			
2	5594	1	143			
2	5595	1	150			
2	5596	1	150			
2	5597	1	150			
2	5598	1	150			
2	5599	1	150			
2	5600	1	150			
2	5601	1	150			
2	5602	1	150			
2	5603	1	159			
2	5604	1	159			
2	5605	1	159			
2	5606	1	159			
2	5607	1	159			
2	5608	1	159			
2	5609	1	159			
2	5610	1	159			
2	5611	1	159			
2	5612	1	169			
2	5613	1	169			
2	5614	1	169			
2	5615	1	169			
2	5616	1	169			
2	5617	1	169			
2	5618	1	169			
2	5619	1	169			
2	5620	1	169			
2	5621	1	179			
2	5622	1	179			
2	5623	1	179			
2	5624	1	179			
2	5625	1	179			
2	5626	1	179			
2	5627	1	179			
2	5628	1	179			
2	5629	1	179			
2	5630	1	179			
2	5631	1	179			
2	5632	1	190			
2	5633	1	190			
2	5634	1	190			
2	5635	1	190			
2	5636	1	190			
2	5637	1	190			
2	5638	1	190			
2	5639	1	190			
2	5640	1	190			
2	5641	1	190			
2	5642	1	200			
2	5643	1	200			
2	5644	1	200			
2	5645	1	200			
2	5646	1	200			
2	5647	1	200			
2	5648	1	200			
2	5649	1	200			
2	5650	1	200			
2	5651	1	200			
2	5652	1	200			
2	5653	1	200			
2	5654	1	213			
2	5655	1	213			
2	5656	1	213			
2	5657	1	213			
2	5658	1	213			
2	5659	1	213			
2	5660	1	213			
2	5661	1	213			
2	5662	1	223			
2	5663	1	223			
2	5664	1	226			
2	5665	1	226			
2	5666	1	226			
2	5667	1	226			
2	5668	1	226			
2	5669	1	226			
2	5670	1	232			
2	5671	1	232			
2	5672	1	232			
2	5673	1	232			
2	5674	1	232			
2	5675	1	232			
2	5676	1	238			
2	5677	1	238			
2	5678	1	238			
2	5679	1	238			
2	5680	1	238			
2	5681	1	238			
2	5682	1	244			
2	5683	1	244			
2	5684	1	244			
2	5685	1	244			
2	5686	1	244			
2	5687	1	244			
2	5688	1	250			
2	5689	1	250			
2	5690	1	250			
2	5691	1	250			
2	5692	1	250			
2	5693	1	250			
2	5694	1	250			
2	5695	1	257			
2	5696	1	257			
2	5697	1	257			
2	5698	1	257			
2	5699	1	257			
2	5700	1	257			
2	5701	1	257			
2	5702	1	264			
2	5703	1	264			
2	5704	1	264			
2	5705	1	264			
2	5706	1	264			
2	5707	1	264			
2	5708	1	270			
2	5709	1	270			
2	5710	1	270			
2	5711	1	270			
2	5712	1	274			
2	5713	1	274			
2	5714	1	274			
2	5715	1	274			
2	5716	1	274			
2	5717	1	274			
2	5718	1	274			
2	5719	1	274			
2	5720	1	283			
2	5721	1	283			
2	5722	1	283			
2	5723	1	283			
2	5724	1	283			
2	5725	1	283			
2	5726	1	283			
2	5727	1	283			
2	5728	1	283			
2	5729	1	283			
2	5730	1	294			
2	5731	1	294			
2	5732	1	294			
2	5733	1	294			
2	5734	1	294			
2	5735	1	294			
2	5736	1	294			
2	5737	1	294			
2	5738	1	303			
2	5739	1	303			
2	5740	1	303			
2	5741	1	303			
2	5742	1	303			
2	5743	1	303			
2	5744	1	303			
2	5745	1	311			
2	5746	1	311			
2	5747	1	311			
2	5748	1	311			
2	5749	1	311			
2	5750	1	317			
2	5751	1	317			
2	5752	1	317			
2	5753	1	317			
2	5754	1	322			
2	5755	1	322			
2	5756	1	322			
2	5757	1	326			
2	5758	1	326			
2	5759	1	330			
2	5760	1	330			
2	5761	1	330			
2	5762	1	330			
2	5763	1	330			
2	5764	1	330			
2	5765	1	330			
2	5766	1	330			
2	5767	1	330			
2	5768	1	330			
2	5769	1	330			
2	5770	1	330			
2	5771	1	330			
2	5772	1	343			
2	5773	1	343			
2	5774	1	343			
2	5775	1	343			
2	5776	1	343			
2	5777	1	343			
2	5778	1	350			
2	5779	1	350			
2	5780	1	665			
2	5781	1	665			
2	5782	1	665			
2	5783	1	665			
2	5784	1	665			
2	5785	1	679			
2	5786	1	679			
2	5787	1	679			
2	5788	1	679			
2	5789	1	686			
2	5790	1	686			
2	5791	1	686			
2	5792	1	686			
2	5793	1	702			
2	5794	1	702			
2	5795	1	702			
2	5796	1	702			
2	5797	1	724			
2	5798	1	724			
2	5799	1	724			
2	5800	1	736			
2	5801	1	736			
2	5802	1	736			
2	5803	1	736			
2	5804	1	749			
2	5805	1	749			
2	5806	1	749			
2	5807	1	749			
2	5808	1	763			
2	5809	1	763			
2	5810	1	763			
2	5811	1	763			
2	5812	1	763			
2	5813	1	769			
2	5814	1	769			
2	5815	1	779			
2	5816	1	779			
2	5817	1	786			
2	5818	1	786			
2	5819	1	786			
2	5820	1	786			
2	5821	1	786			
2	5822	1	786			
2	5823	1	794			
2	5824	1	794			
2	5825	1	794			
2	5826	1	803			
2	5827	1	803			
2	5828	1	803			
2	5829	1	803			
2	5830	1	803			
2	5831	1	803			
2	5832	1	803			
2	5833	1	803			
2	5834	1	803			
2	5835	1	803			
2	5836	1	803			
2	5837	1	803			
2	5838	1	803			
2	5839	1	803			
2	5840	1	803			
2	5841	1	803			
2	5842	1	825			
2	5843	1	825			
2	5844	1	825			
2	5845	1	825			
2	5846	1	825			
2	5847	1	825			
2	5848	1	825			
2	5849	1	825			
2	5850	1	825			
2	5851	1	825			
2	5852	1	825			
2	5853	1	825			
2	5854	1	825			
2	5855	1	825			
2	5856	1	825			
2	5857	1	825			
2	5858	1	825			
2	5859	1	825			
2	5860	1	825			
2	5861	1	825			
2	5862	1	829			
2	5863	1	829			
2	5864	1	832			
2	5865	1	832			
2	5866	1	832			
2	5867	1	832			
2	5868	1	839			
2	5869	1	839			
2	5870	1	839			
2	5871	1	839			
2	5872	1	842			
2	5873	1	842			
2	5874	1	848			
2	5875	1	848			
2	5876	1	854			
2	5877	1	854			
2	5878	1	854			
2	5879	1	861			
2	5880	1	861			
2	5881	1	867			
2	5882	1	867			
2	5883	1	870			
2	5884	1	870			
2	5885	1	870			
2	5886	1	883			
2	5887	1	883			
2	5888	1	892			
2	5889	1	892			
2	5890	1	892			
2	5891	1	896			
2	5892	1	896			
2	5893	1	896			
2	5894	1	896			
2	5895	1	896			
2	5896	1	896			
2	5897	1	896			
2	5898	1	896			
2	5899	1	896			
2	5900	1	896			
2	5901	1	896			
2	5902	1	896			
2	5903	1	896			
2	5904	1	896			
2	5905	1	896			
2	5906	1	896			
2	5907	1	920			
2	5908	1	920			
2	5909	1	1117			
2	5910	1	1117			
2	5911	1	1117			
2	5912	1	1117			
2	5913	1	1117			
2	5914	1	1117			
2	5915	1	1117			
2	5916	1	1117			
2	5917	1	1117			
2	5918	1	1117			
2	5919	1	1117			
2	5920	1	1117			
2	5921	1	1117			
2	5922	1	1117			
2	5923	1	1117			
2	5924	1	1117			
2	5925	1	1197			
2	5926	1	1197			
2	5927	1	1197			
2	5928	1	1197			
2	5929	1	1202			
2	5930	1	1202			
2	5931	1	1202			
2	5932	1	1202			
2	5933	1	1202			
2	5934	1	1202			
2	5935	1	1202			
2	5936	1	1202			
2	5937	1	1202			
2	5938	1	1202			
2	5939	1	1202			
2	5940	1	1202			
2	5941	1	1202			
2	5942	1	1202			
2	5943	1	1202			
2	5944	1	1202			
2	5945	1	1219			
2	5946	1	1219			
2	5947	1	1219			
2	5948	1	1219			
2	5949	1	1264			
2	5950	1	1264			
2	5951	1	1306			
2	5952	1	1306			
2	5953	1	1306			
2	5954	1	1306			
2	5955	1	1306			
2	5956	1	1306			
2	5957	1	1306			
2	5958	1	1306			
2	5959	1	1315			
2	5960	1	1315			
2	5961	1	1315			
2	5962	1	1315			
2	5963	1	1315			
2	5964	1	1315			
2	5965	1	1322			
2	5966	1	1322			
2	5967	1	1325			
2	5968	1	1325			
2	5969	1	1328			
2	5970	1	1328			
2	5971	1	1331			
2	5972	1	1331			
2	5973	1	1340			
2	5974	1	1340			
2	5975	1	1353			
2	5976	1	1353			
2	5977	1	1353			
2	5978	1	1353			
2	5979	1	1358			
2	5980	1	1358			
2	5981	1	1358			
2	5982	1	1358			
2	5983	1	1366			
2	5984	1	1366			
2	5985	1	1409			
2	5986	1	1409			
2	5987	1	1409			
2	5988	1	1409			
2	5989	1	1409			
2	5990	1	1409			
2	5991	1	1409			
2	5992	1	1409			
2	5993	1	1409			
2	5994	1	1409			
2	5995	1	1409			
2	5996	1	1409			
2	5997	1	1409			
2	5998	1	1409			
2	5999	1	1409			
2	6000	1	1409			
2	6001	1	1452			
2	6002	1	1452			
2	6003	1	1452			
2	6004	1	1452			
2	6005	1	1452			
2	6006	1	1452			
2	6007	1	1461			
2	6008	1	1461			
2	6009	1	1464			
2	6010	1	1464			
2	6011	1	1464			
2	6012	1	1520			
2	6013	1	1520			
2	6014	1	1520			
2	6015	1	1562			
2	6016	1	1562			
2	6017	1	1562			
2	6018	1	1562			
2	6019	1	1562			
2	6020	1	1562			
2	6021	1	1562			
2	6022	1	1562			
2	6023	1	1562			
2	6024	1	1562			
2	6025	1	1562			
2	6026	1	1562			
2	6027	1	1562			
2	6028	1	1562			
2	6029	1	1562			
2	6030	1	1562			
2	6031	1	1667			
2	6032	1	1667			
2	6033	1	1667			
2	6034	1	1667			
2	6035	1	1667			
2	6036	1	1670			
2	6037	1	1670			
2	6038	1	1670			
2	6039	1	1670			
2	6040	1	1670			
2	6041	1	1715			
2	6042	1	1715			
2	6043	1	1715			
2	6044	1	1715			
2	6045	1	1718			
2	6046	1	1718			
2	6047	1	1718			
2	6048	1	1718			
2	6049	1	1722			
2	6050	1	1722			
2	6051	1	1738			
2	6052	1	1738			
2	6053	1	1738			
2	6054	1	1738			
2	6055	1	1738			
2	6056	1	1738			
2	6057	1	1738			
2	6058	1	1738			
2	6059	1	1747			
2	6060	1	1747			
2	6061	1	1747			
2	6062	1	1747			
2	6063	1	1747			
2	6064	1	1747			
2	6065	1	1747			
2	6066	1	1747			
2	6067	1	1756			
2	6068	1	1756			
2	6069	1	1756			
2	6070	1	1756			
2	6071	1	1761			
2	6072	1	1761			
2	6073	1	1761			
2	6074	1	1761			
2	6075	1	1761			
2	6076	1	1761			
2	6077	1	1761			
2	6078	1	1761			
2	6079	1	1761			
2	6080	1	1761			
2	6081	1	1761			
2	6082	1	1761			
2	6083	1	1761			
2	6084	1	1761			
2	6085	1	1761			
2	6086	1	1761			
2	6087	1	1761			
2	6088	1	1761			
2	6089	1	1803			
2	6090	1	1803			
2	6091	1	1806			
2	6092	1	1806			
2	6093	1	1809			
2	6094	1	1809			
2	6095	1	1812			
2	6096	1	1812			
2	6097	1	1815			
2	6098	1	1815			
2	6099	1	1818			
2	6100	1	1818			
2	6101	1	1821			
2	6102	1	1821			
2	6103	1	1821			
2	6104	1	1821			
2	6105	1	1821			
2	6106	1	1821			
2	6107	1	1821			
2	6108	1	1821			
2	6109	1	1821			
2	6110	1	1821			
2	6111	1	1821			
2	6112	1	1821			
2	6113	1	1821			
2	6114	1	1821			
2	6115	1	1821			
2	6116	1	1821			
2	6117	1	1824			
2	6118	1	1824			
2	6119	1	1824			
2	6120	1	1824			
2	6121	1	1824			
2	6122	1	1824			
2	6123	1	1824			
2	6124	1	1824			
2	6125	1	1833			
2	6126	1	1833			
2	6127	1	1833			
2	6128	1	1833			
2	6129	1	1833			
2	6130	1	1833			
2	6131	1	1833			
2	6132	1	1833			
2	6133	1	1870			
2	6134	1	1870			
2	6135	1	1875			
2	6136	1	1875			
2	6137	1	1880			
2	6138	1	1880			
2	6139	1	1885			
2	6140	1	1885			
2	6141	1	1890			
2	6142	1	1890			
2	6143	1	1895			
2	6144	1	1895			
2	6145	1	1900			
2	6146	1	1900			
2	6147	1	1905			
2	6148	1	1905			
2	6149	1	1909			
2	6150	1	1909			
2	6151	1	1913			
2	6152	1	1913			
2	6153	1	1913			
2	6154	1	1917			
2	6155	1	1917			
2	6156	1	1917			
2	6157	1	1917			
2	6158	1	1917			
2	6159	1	1922			
2	6160	1	1922			
2	6161	1	1922			
2	6162	1	1926			
2	6163	1	1926			
2	6164	1	1926			
2	6165	1	1933			
2	6166	1	1933			
2	6167	1	1936			
2	6168	1	1936			
2	6169	1	1983			
2	6170	1	1983			
2	6171	1	2043			
2	6172	1	2043			
2	6173	1	2043			
2	6174	1	2043			
2	6175	1	2043			
2	6176	1	2043			
2	6177	1	2043			
2	6178	1	2043			
2	6179	1	2057			
2	6180	1	2057			
2	6181	1	2057			
2	6182	1	2057			
2	6183	1	2057			
2	6184	1	2057			
2	6185	1	2057			
2	6186	1	2057			
2	6187	1	2068			
2	6188	1	2068			
2	6189	1	2073			
2	6190	1	2073			
2	6191	1	2078			
2	6192	1	2078			
2	6193	1	2083			
2	6194	1	2083			
2	6195	1	2088			
2	6196	1	2088			
2	6197	1	2093			
2	6198	1	2093			
2	6199	1	2098			
2	6200	1	2098			
2	6201	1	2103			
2	6202	1	2103			
2	6203	1	2185			
2	6204	1	2185			
2	6205	1	2185			
2	6206	1	2185			
2	6207	1	2185			
2	6208	1	2185			
2	6209	1	2185			
2	6210	1	2185			
2	6211	1	2185			
2	6212	1	2185			
2	6213	1	2185			
2	6214	1	2185			
2	6215	1	2185			
2	6216	1	2185			
2	6217	1	2185			
2	6218	1	2185			
2	6219	1	2188			
2	6220	1	2188			
2	6221	1	2188			
2	6222	1	2188			
2	6223	1	2188			
2	6224	1	2188			
2	6225	1	2188			
2	6226	1	2188			
2	6227	1	2188			
2	6228	1	2188			
2	6229	1	2188			
2	6230	1	2188			
2	6231	1	2188			
2	6232	1	2188			
2	6233	1	2188			
2	6234	1	2188			
2	6235	1	2191			
2	6236	1	2191			
2	6237	1	2191			
2	6238	1	2191			
2	6239	1	2191			
2	6240	1	2191			
2	6241	1	2191			
2	6242	1	2191			
2	6243	1	2191			
2	6244	1	2191			
2	6245	1	2191			
2	6246	1	2191			
2	6247	1	2191			
2	6248	1	2191			
2	6249	1	2191			
2	6250	1	2191			
2	6251	1	2194			
2	6252	1	2194			
2	6253	1	2194			
2	6254	1	2194			
2	6255	1	2194			
2	6256	1	2194			
2	6257	1	2194			
2	6258	1	2194			
2	6259	1	2194			
2	6260	1	2194			
2	6261	1	2194			
2	6262	1	2194			
2	6263	1	2194			
2	6264	1	2194			
2	6265	1	2194			
2	6266	1	2194			
2	6267	1	2197			
2	6268	1	2197			
2	6269	1	2197			
2	6270	1	2197			
2	6271	1	2197			
2	6272	1	2197			
2	6273	1	2197			
2	6274	1	2197			
2	6275	1	2197			
2	6276	1	2197			
2	6277	1	2197			
2	6278	1	2197			
2	6279	1	2197			
2	6280	1	2197			
2	6281	1	2197			
2	6282	1	2197			
2	6283	1	2200			
2	6284	1	2200			
2	6285	1	2200			
2	6286	1	2200			
2	6287	1	2200			
2	6288	1	2200			
2	6289	1	2200			
2	6290	1	2200			
2	6291	1	2200			
2	6292	1	2200			
2	6293	1	2200			
2	6294	1	2200			
2	6295	1	2200			
2	6296	1	2200			
2	6297	1	2200			
2	6298	1	2200			
2	6299	1	2203			
2	6300	1	2203			
2	6301	1	2203			
2	6302	1	2203			
2	6303	1	2203			
2	6304	1	2203			
2	6305	1	2203			
2	6306	1	2203			
2	6307	1	2203			
2	6308	1	2203			
2	6309	1	2203			
2	6310	1	2203			
2	6311	1	2203			
2	6312	1	2203			
2	6313	1	2203			
2	6314	1	2203			
2	6315	1	2206			
2	6316	1	2206			
2	6317	1	2206			
2	6318	1	2206			
2	6319	1	2206			
2	6320	1	2206			
2	6321	1	2206			
2	6322	1	2206			
2	6323	1	2206			
2	6324	1	2206			
2	6325	1	2206			
2	6326	1	2206			
2	6327	1	2206			
2	6328	1	2206			
2	6329	1	2206			
2	6330	1	2206			
2	6331	1	2270			
2	6332	1	2270			
2	6333	1	2277			
2	6334	1	2277			
2	6335	1	2282			
2	6336	1	2282			
2	6337	1	2287			
2	6338	1	2287			
2	6339	1	2294			
2	6340	1	2294			
2	6341	1	2299			
2	6342	1	2299			
2	6343	1	2307			
2	6344	1	2307			
2	6345	1	2310			
2	6346	1	2310			
2	6347	1	2325			
2	6348	1	2325			
2	6349	1	2328			
2	6350	1	2328			
2	6351	1	2331			
2	6352	1	2331			
2	6353	1	2334			
2	6354	1	2334			
2	6355	1	2376			
2	6356	1	2376			
2	6357	1	2379			
2	6358	1	2379			
2	6359	1	2471			
2	6360	1	2471			
2	6361	1	2471			
2	6362	1	2471			
2	6363	1	2471			
2	6364	1	2483			
2	6365	1	2483			
2	6366	1	2648			
2	6367	1	2648			
2	6368	1	2648			
2	6369	1	2652			
2	6370	1	2652			
2	6371	1	2652			
2	6372	1	2656			
2	6373	1	2656			
2	6374	1	2656			
2	6375	1	2659			
2	6376	1	2659			
2	6377	1	2659			
2	6378	1	2662			
2	6379	1	2662			
2	6380	1	2662			
2	6381	1	2666			
2	6382	1	2666			
2	6383	1	2666			
2	6384	1	2670			
2	6385	1	2670			
2	6386	1	2670			
2	6387	1	2673			
2	6388	1	2673			
2	6389	1	2673			
2	6390	1	2677			
2	6391	1	2677			
2	6392	1	2677			
2	6393	1	2681			
2	6394	1	2681			
2	6395	1	2681			
2	6396	1	2684			
2	6397	1	2684			
2	6398	1	2684			
2	6399	1	2688			
2	6400	1	2688			
2	6401	1	2688			
2	6402	1	2692			
2	6403	1	2692			
2	6404	1	2692			
2	6405	1	2692			
2	6406	1	2692			
2	6407	1	2697			
2	6408	1	2697			
2	6409	1	2697			
2	6410	1	2697			
2	6411	1	2697			
2	6412	1	2702			
2	6413	1	2702			
2	6414	1	2702			
2	6415	1	2706			
2	6416	1	2706			
2	6417	1	2706			
2	6418	1	2710			
2	6419	1	2710			
2	6420	1	2710			
2	6421	1	2710			
2	6422	1	2710			
2	6423	1	2715			
2	6424	1	2715			
2	6425	1	2715			
2	6426	1	2719			
2	6427	1	2719			
2	6428	1	2719			
2	6429	1	2723			
2	6430	1	2723			
2	6431	1	2723			
2	6432	1	2723			
2	6433	1	2723			
2	6434	1	2758			
2	6435	1	2758			
2	6436	1	2761			
2	6437	1	2761			
2	6438	1	2764			
2	6439	1	2764			
2	6440	1	2967			
2	6441	1	2967			
2	6442	1	2967			
2	6443	1	2967			
2	6444	1	2973			
2	6445	1	2973			
2	6446	1	2973			
2	6447	1	2973			
2	6448	1	2973			
2	6449	1	2977			
2	6450	1	2977			
2	6451	1	2977			
2	6452	1	2977			
2	6453	1	2977			
2	6454	1	3115			
2	6455	1	3115			
2	6456	1	3119			
2	6457	1	3119			
2	6458	1	3125			
2	6459	1	3125			
2	6460	1	3131			
2	6461	1	3131			
2	6462	1	3138			
2	6463	1	3138			
2	6464	1	3145			
2	6465	1	3145			
2	6466	1	3149			
2	6467	1	3149			
2	6468	1	3155			
2	6469	1	3155			
2	6470	1	3161			
2	6471	1	3161			
2	6472	1	3168			
2	6473	1	3168			
2	6474	1	3172			
2	6475	1	3172			
2	6476	1	3172			
2	6477	1	3172			
2	6478	1	3175			
2	6479	1	3175			
2	6480	1	3175			
2	6481	1	3175			
2	6482	1	3178			
2	6483	1	3178			
2	6484	1	3178			
2	6485	1	3178			
2	6486	1	3181			
2	6487	1	3181			
2	6488	1	3181			
2	6489	1	3181			
2	6490	1	3184			
2	6491	1	3184			
2	6492	1	3184			
2	6493	1	3184			
2	6494	1	3187			
2	6495	1	3187			
2	6496	1	3187			
2	6497	1	3187			
2	6498	1	3407			
2	6499	1	3407			
2	6500	1	3410			
2	6501	1	3410			
2	6502	1	3415			
2	6503	1	3415			
2	6504	1	3415			
2	6505	1	3419			
2	6506	1	3419			
2	6507	1	3419			
2	6508	1	3423			
2	6509	1	3423			
2	6510	1	3426			
2	6511	1	3426			
2	6512	1	3431			
2	6513	1	3431			
2	6514	1	3434			
2	6515	1	3434			
2	6516	1	3439			
2	6517	1	3439			
2	6518	1	3442			
2	6519	1	3442			
2	6520	1	3447			
2	6521	1	3447			
2	6522	1	3447			
2	6523	1	3451			
2	6524	1	3451			
2	6525	1	3451			
2	6526	1	3455			
2	6527	1	3455			
2	6528	1	3458			
2	6529	1	3458			
2	6530	1	3463			
2	6531	1	3463			
2	6532	1	3466			
2	6533	1	3466			
2	6534	1	3645			
2	6535	1	3645			
2	6536	1	3648			
2	6537	1	3648			
2	6538	1	3654			
2	6539	1	3654			
2	6540	1	3658			
2	6541	1	3658			
2	6542	1	3664			
2	6543	1	3664			
2	6544	1	3667			
2	6545	1	3667			
2	6546	1	3673			
2	6547	1	3673			
2	6548	1	3677			
2	6549	1	3677			
2	6550	1	3682			
2	6551	1	3682			
2	6552	1	3682			
2	6553	1	3682			
2	6554	1	3690			
2	6555	1	3690			
2	6556	1	3690			
2	6557	1	3690			
2	6558	1	3721			
2	6559	1	3721			
2	6560	1	3721			
2	6561	1	3721			
2	6562	1	3721			
2	6563	1	3721			
2	6564	1	3721			
2	6565	1	3721			
2	6566	1	3734			
2	6567	1	3734			
2	6568	1	3734			
2	6569	1	3734			
2	6570	1	3734			
2	6571	1	3734			
2	6572	1	3740			
2	6573	1	3740			
2	6574	1	3740			
2	6575	1	3740			
2	6576	1	3740			
2	6577	1	3743			
2	6578	1	3743			
2	6579	1	3743			
2	6580	1	3743			
2	6581	1	3743			
2	6582	1	3743			
2	6583	1	3743			
2	6584	1	3743			
2	6585	1	3756			
2	6586	1	3756			
2	6587	1	3756			
2	6588	1	3756			
2	6589	1	3756			
2	6590	1	3756			
2	6591	1	3762			
2	6592	1	3762			
2	6593	1	3762			
2	6594	1	3762			
2	6595	1	3762			
2	6596	1	3786			
2	6597	1	3786			
2	6598	1	3800			
2	6599	1	3800			
2	6600	1	3809			
2	6601	1	3809			
2	6602	1	3812			
2	6603	1	3812			
2	6604	1	3812			
2	6605	1	3815			
2	6606	1	3815			
2	6607	1	3818			
2	6608	1	3818			
2	6609	1	3818			
2	6610	1	3818			
2	6611	1	3838			
2	6612	1	3838			
2	6613	1	3838			
2	6614	1	3838			
2	6615	1	3838			
2	6616	1	3838			
2	6617	1	3838			
2	6618	1	3845			
2	6619	1	3845			
2	6620	1	3845			
2	6621	1	3845			
2	6622	1	3845			
2	6623	1	3845			
2	6624	1	3845			
2	6625	1	3926			
2	6626	1	3926			
2	6627	1	3926			
2	6628	1	3926			
2	6629	1	3932			
2	6630	1	3932			
2	6631	1	3992			
2	6632	1	3992			
2	6633	1	3996			
2	6634	1	3996			
2	6635	1	4091			
2	6636	1	4091			
2	6637	1	4091			
2	6638	1	4091			
2	6639	1	4091			
2	6640	1	4091			
2	6641	1	4091			
2	6642	1	4091			
2	6643	1	4091			
2	6644	1	4094			
2	6645	1	4094			
2	6646	1	4094			
2	6647	1	4094			
2	6648	1	4094			
2	6649	1	4094			
2	6650	1	4116			
2	6651	1	4116			
2	6652	1	4116			
2	6653	1	4116			
2	6654	1	4116			
2	6655	1	4116			
2	6656	1	4116			
2	6657	1	4116			
2	6658	1	4119			
2	6659	1	4119			
2	6660	1	4119			
2	6661	1	4119			
2	6662	1	4119			
2	6663	1	4119			
2	6664	1	4119			
2	6665	1	4119			
2	6666	1	4123			
2	6667	1	4123			
2	6668	1	4123			
2	6669	1	4123			
2	6670	1	4123			
2	6671	1	4128			
2	6672	1	4128			
2	6673	1	4128			
2	6674	1	4128			
2	6675	1	4128			
2	6676	1	4128			
2	6677	1	4139			
2	6678	1	4139			
2	6679	1	4142			
2	6680	1	4142			
2	6681	1	4186			
2	6682	1	4186			
2	6683	1	4197			
2	6684	1	4197			
2	6685	1	4197			
2	6686	1	4197			
2	6687	1	4197			
2	6688	1	4197			
2	6689	1	4218			
2	6690	1	4218			
2	6691	1	4218			
2	6692	1	4218			
2	6693	1	4218			
2	6694	1	4242			
2	6695	1	4242			
2	6696	1	4242			
2	6697	1	4242			
2	6698	1	4284			
2	6699	1	4284			
2	6700	1	4284			
2	6701	1	4287			
2	6702	1	4287			
2	6703	1	4287			
2	6704	1	4287			
2	6705	1	4287			
2	6706	1	4310			
2	6707	1	4310			
2	6708	1	4310			
2	6709	1	4310			
2	6710	1	4310			
2	6711	1	4319			
2	6712	1	4319			
2	6713	1	4331			
2	6714	1	4331			
2	6715	1	4335			
2	6716	1	4335			
2	6717	1	4338			
2	6718	1	4338			
2	6719	1	4341			
2	6720	1	4341			
2	6721	1	4344			
2	6722	1	4344			
2	6723	1	4347			
2	6724	1	4347			
2	6725	1	4350			
2	6726	1	4350			
2	6727	1	4371			
2	6728	1	4371			
2	6729	1	4387			
2	6730	1	4387			
2	6731	1	4387			
2	6732	1	4387			
2	6733	1	4390			
2	6734	1	4390			
2	6735	1	4390			
2	6736	1	4390			
2	6737	1	4416			
2	6738	1	4416			
2	6739	1	4421			
2	6740	1	4421			
2	6741	1	4427			
2	6742	1	4427			
2	6743	1	4435			
2	6744	1	4435			
2	6745	1	4443			
2	6746	1	4443			
2	6747	1	4443			
2	6748	1	4458			
2	6749	1	4458			
2	6750	1	4458			
2	6751	1	4458			
2	6752	1	4468			
2	6753	1	4468			
2	6754	1	4468			
2	6755	1	4468			
2	6756	1	4468			
2	6757	1	4472			
2	6758	1	4472			
2	6759	1	4475			
2	6760	1	4475			
2	6761	1	4493			
2	6762	1	4493			
2	6763	1	4498			
2	6764	1	4498			
2	6765	1	4503			
2	6766	1	4503			
2	6767	1	4503			
2	6768	1	4503			
2	6769	1	4549			
2	6770	1	4549			
2	6771	1	4549			
2	6772	1	4549			
2	6773	1	4559			
2	6774	1	4559			
2	6775	1	4576			
2	6776	1	4576			
2	6777	1	4593			
2	6778	1	4593			
2	6779	1	4593			
2	6780	1	4593			
2	6781	1	4599			
2	6782	1	4599			
2	6783	1	4599			
2	6784	1	4599			
2	6785	1	4619			
2	6786	1	4619			
2	6787	1	4623			
2	6788	1	4623			
2	6789	1	4644			
2	6790	1	4644			
2	6791	1	4644			
2	6792	1	4644			
2	6793	1	4644			
2	6794	1	4647			
2	6795	1	4647			
2	6796	1	4650			
2	6797	1	4650			
2	6798	1	4711			
2	6799	1	4711			
2	6800	1	4717			
2	6801	1	4717			
2	6802	1	4717			
2	6803	1	4727			
2	6804	1	4727			
2	6805	1	4727			
2	6806	1	4730			
2	6807	1	4730			
2	6808	1	4740			
2	6809	1	4740			
2	6810	1	4740			
2	6811	1	4740			
2	6812	1	4743			
2	6813	1	4743			
2	6814	1	4743			
2	6815	1	4743			
2	6816	1	4757			
2	6817	1	4757			
2	6818	1	4757			
2	6819	1	4757			
2	6820	1	4769			
2	6821	1	4769			
2	6822	1	4772			
2	6823	1	4772			
2	6824	1	4775			
2	6825	1	4775			
2	6826	1	4794			
2	6827	1	4794			
2	6828	1	4797			
2	6829	1	4797			
2	6830	1	4800			
2	6831	1	4800			
2	6832	1	4808			
2	6833	1	4808			
2	6834	1	4818			
2	6835	1	4818			
2	6836	1	4818			
2	6837	1	4823			
2	6838	1	4823			
2	6839	1	4831			
2	6840	1	4831			
2	6841	1	4838			
2	6842	1	4838			
2	6843	1	4876			
2	6844	1	4876			
2	6845	1	4876			
2	6846	1	4876			
2	6847	1	4876			
2	6848	1	4880			
2	6849	1	4880			
2	6850	1	4889			
2	6851	1	4889			
2	6852	1	4907			
2	6853	1	4907			
2	6854	1	4913			
2	6855	1	4913			
2	6856	1	4916			
2	6857	1	4916			
2	6858	1	4921			
2	6859	1	4921			
2	6860	1	4946			
2	6861	1	4946			
2	6862	1	4954			
2	6863	1	4954			
2	6864	1	4957			
2	6865	1	4957			
2	6866	1	4973			
2	6867	1	4973			
2	6868	1	4985			
2	6869	1	4985			
2	6870	1	4988			
2	6871	1	4988			
2	6872	1	4988			
2	6873	1	4991			
2	6874	1	4991			
2	6875	1	4996			
2	6876	1	4996			
2	6877	1	4996			
2	6878	1	4999			
2	6879	1	4999			
2	6880	1	5010			
2	6881	1	5010			
2	6882	1	5013			
2	6883	1	5013			
2	6884	1	5018			
2	6885	1	5018			
2	6886	1	5018			
2	6887	1	5021			
2	6888	1	5021			
2	6889	1	5030			
2	6890	1	5030			
2	6891	1	5050			
2	6892	1	5050			
2	6893	1	5050			
2	6894	1	5050			
2	6895	1	5050			
2	6896	1	5055			
2	6897	1	5055			
2	6898	1	5058			
2	6899	1	5058			
2	6900	1	5058			
2	6901	1	5058			
2	6902	1	5058			
2	6903	1	5061			
2	6904	1	5061			
2	6905	1	5066			
2	6906	1	5066			
2	6907	1	5080			
2	6908	1	5080			
2	6909	1	5080			
2	6910	1	5080			
2	6911	1	5080			
2	6912	1	5085			
2	6913	1	5085			
2	6914	1	5114			
2	6915	1	5114			
2	6916	1	5114			
2	6917	1	5114			
2	6918	1	5122			
2	6919	1	5122			
2	6920	1	5122			
2	6921	1	5122			
2	6922	1	5128			
2	6923	1	5128			
2	6924	1	5128			
2	6925	1	5128			
2	6926	1	5133			
2	6927	1	5133			
2	6928	1	5145			
2	6929	1	5145			
2	6930	1	5145			
2	6931	1	5145			
2	6932	1	5228			
2	6933	1	5228			
2	6934	1	5236			
2	6935	1	5236			
2	6936	1	5236			
2	6937	1	5236			
2	6938	1	5250			
2	6939	1	5250			
2	6940	1	5254			
2	6941	1	5254			
2	6942	1	5258			
2	6943	1	5258			
2	6944	1	5258			
2	6945	1	5258			
2	6946	1	5266			
2	6947	1	5266			
2	6948	1	5279			
2	6949	1	5279			
2	6950	1	5279			
2	6951	1	5279			
2	6952	1	5298			
2	6953	1	5298			
2	6954	1	5298			
2	6955	1	5298			
2	6956	1	5309			
2	6957	1	5309			
2	6958	1	5309			
2	6959	1	5309			
