1 1 0 2 0
1 4 0 2 0
1 7 0 2 0
1 10 0 2 0
1 13 0 2 0
1 16 0 2 0
1 19 0 2 0
1 22 0 2 0
1 25 0 2 0
1 28 0 2 0
1 31 0 2 0
1 34 0 2 0
1 37 0 2 0
1 40 0 2 0
1 43 0 2 0
1 46 0 2 0
1 49 0 3 0
1 53 0 2 0
1 56 0 3 0
1 60 0 2 0
1 63 0 2 0
1 66 0 2 0
1 69 0 2 0
1 72 0 3 0
1 76 0 2 0
1 79 0 2 0
1 82 0 2 0
1 85 0 2 0
1 88 0 2 0
1 91 0 2 0
1 94 0 4 0
1 99 0 4 0
1 104 0 7 0
0 190 5 3 1 2
0 194 5 2 1 5
0 197 5 3 1 8
0 201 5 4 1 11
0 206 5 2 1 14
0 209 5 2 1 17
0 212 5 3 1 20
0 216 5 3 1 23
0 220 5 4 1 26
0 225 5 3 1 29
0 229 5 2 1 32
0 232 5 2 1 35
0 235 5 3 1 38
0 239 5 3 1 41
0 243 5 3 1 44
0 247 5 3 1 47
0 251 6 1 2 64 89
0 252 6 1 2 67 92
0 253 5 2 1 73
0 256 5 1 1 74
0 257 1 2 1 70
0 260 1 2 1 71
0 263 5 2 1 77
0 266 5 2 1 80
0 269 5 2 1 83
0 272 5 2 1 86
0 275 5 1 1 105
0 276 5 1 1 106
0 277 5 2 1 90
0 280 5 2 1 93
0 283 1 6 1 95
0 290 5 6 1 96
0 297 1 2 1 97
0 300 5 2 1 98
0 303 1 2 1 100
0 306 5 6 1 101
0 313 5 2 1 102
0 316 1 2 1 107
0 319 5 6 1 108
0 326 1 4 1 109
0 331 1 6 1 110
0 338 5 4 1 111
0 343 1 2 1 3
0 346 1 2 1 6
0 349 1 2 1 9
0 352 1 2 1 12
0 355 1 2 1 15
0 358 1 2 1 18
0 361 1 2 1 21
0 364 1 2 1 24
0 367 1 2 1 27
0 370 1 2 1 30
0 373 1 2 1 33
0 376 1 2 1 36
0 379 1 2 1 39
0 382 1 2 1 42
0 385 1 2 1 45
0 388 1 2 1 48
0 534 5 1 1 236
0 535 5 1 1 238
0 536 5 1 1 241
0 537 5 1 1 244
0 538 5 1 1 246
0 539 5 1 1 249
0 540 5 1 1 254
0 541 5 1 1 258
0 542 5 1 1 261
0 543 5 1 1 264
0 544 5 1 1 267
0 545 5 1 1 270
0 546 5 1 1 273
0 547 5 1 1 278
0 548 5 1 1 281
0 549 5 1 1 284
0 550 6 1 2 195 222
0 551 6 1 2 196 223
0 552 6 1 2 198 224
0 553 6 1 2 199 226
0 554 6 1 2 200 227
0 555 6 1 2 202 228
0 556 1 2 1 112
0 559 1 2 1 115
0 562 1 2 1 124
0 565 1 2 1 126
0 568 1 2 1 138
0 571 1 2 1 151
0 574 7 2 2 65 208
0 577 1 2 1 134
0 580 1 2 1 141
0 583 1 2 1 143
0 586 7 2 2 68 210
0 589 1 2 1 148
0 592 7 2 3 50 157 211
0 595 1 2 1 154
0 598 1 2 1 149
0 601 6 1 2 217 171
0 602 6 1 2 218 173
0 603 6 4 2 161 75
0 608 6 3 2 162 189
0 612 6 3 2 256 191
0 616 1 2 1 120
0 619 1 2 1 131
0 622 1 2 1 135
0 625 1 2 1 150
0 628 1 2 1 113
0 631 1 2 1 114
0 634 1 2 1 116
0 637 1 2 1 142
0 640 1 2 1 117
0 643 7 2 3 57 159 213
0 646 1 2 1 144
0 649 1 2 1 121
0 652 1 2 1 145
0 655 7 2 3 61 160 214
0 658 1 2 1 163
0 661 1 2 1 164
0 664 1 2 1 165
0 667 1 2 1 166
0 670 1 2 1 167
0 673 1 2 1 168
0 676 1 2 1 169
0 679 1 2 1 170
0 682 7 2 2 251 205
0 685 7 2 2 252 207
0 688 1 2 1 118
0 691 1 2 1 119
0 694 1 2 1 128
0 697 1 2 1 129
0 700 1 2 1 155
0 703 1 2 1 156
0 706 1 2 1 146
0 709 1 2 1 147
0 712 1 2 1 122
0 715 1 2 1 123
0 718 1 2 1 125
0 721 1 2 1 132
0 724 7 2 3 54 158 215
0 727 1 2 1 152
0 730 1 2 1 136
0 733 1 2 1 137
0 736 1 2 1 127
0 739 1 2 1 133
0 742 1 2 1 139
0 745 1 2 1 153
0 748 1 2 1 130
0 751 1 2 1 140
0 886 5 1 1 397
0 887 5 1 1 399
0 888 5 1 1 336
0 889 5 1 1 339
0 890 5 1 1 341
0 891 5 1 1 344
0 892 5 1 1 350
0 893 5 1 1 362
0 894 5 1 1 368
0 895 5 1 1 371
0 896 5 1 1 374
0 897 7 1 2 51 333
0 898 7 1 2 58 329
0 899 6 3 2 55 334
0 903 6 3 2 62 330
0 907 6 2 2 52 335
0 910 6 2 2 59 332
0 913 5 1 1 380
0 914 5 1 1 377
0 915 5 1 1 386
0 916 5 1 1 383
0 917 5 1 1 391
0 918 5 1 1 389
0 919 5 1 1 395
0 920 5 1 1 393
0 921 6 1 4 172 187 219 324
0 922 6 1 4 174 188 221 325
0 923 6 2 3 192 230 327
0 926 7 8 3 193 231 328
0 935 1 2 1 286
0 938 5 1 1 401
0 939 1 2 1 287
0 942 5 1 1 403
0 943 1 2 1 291
0 946 5 1 1 405
0 947 1 2 1 292
0 950 5 1 1 407
0 951 1 2 1 295
0 954 5 1 1 409
0 955 1 2 1 296
0 958 5 1 1 411
0 959 1 2 1 301
0 962 1 2 1 302
0 965 1 2 1 307
0 968 5 1 1 413
0 969 1 2 1 308
0 972 5 1 1 415
0 973 1 2 1 311
0 976 5 1 1 417
0 977 1 2 1 312
0 980 5 1 1 419
0 981 1 2 1 317
0 984 5 1 1 347
0 985 1 2 1 318
0 988 5 1 1 421
0 989 5 1 1 423
0 990 5 1 1 353
0 991 5 1 1 425
0 992 5 1 1 427
0 993 5 1 1 356
0 994 1 2 1 320
0 997 5 1 1 429
0 998 1 2 1 321
0 1001 5 1 1 431
0 1002 5 1 1 433
0 1003 5 1 1 435
0 1004 5 1 1 359
0 1005 5 1 1 437
0 1006 5 1 1 439
0 1007 5 1 1 365
0 1008 5 1 1 441
0 1009 5 1 1 443
0 1010 1 2 1 288
0 1013 1 2 1 289
0 1016 1 2 1 293
0 1019 1 2 1 294
0 1022 1 2 1 298
0 1025 1 2 1 299
0 1028 1 2 1 304
0 1031 1 2 1 305
0 1034 1 2 1 309
0 1037 1 2 1 310
0 1040 1 2 1 314
0 1043 1 2 1 315
0 1046 1 2 1 322
0 1049 1 2 1 323
0 1054 6 1 2 340 888
0 1055 6 1 2 337 889
0 1063 6 1 2 345 890
0 1064 6 1 2 342 891
0 1067 6 1 2 375 895
0 1068 6 1 2 372 896
0 1119 6 1 2 424 988
0 1120 6 1 2 422 989
0 1121 6 1 2 428 991
0 1122 6 1 2 426 992
0 1128 6 1 2 436 1002
0 1129 6 1 2 434 1003
0 1130 6 1 2 440 1005
0 1131 6 1 2 438 1006
0 1132 6 1 2 444 1008
0 1133 6 1 2 442 1009
0 1148 5 1 1 467
0 1149 5 1 1 465
0 1150 6 1 2 1054 1055
0 1151 5 1 1 469
0 1152 5 1 1 471
0 1153 5 1 1 475
0 1154 5 1 1 473
0 1155 5 1 1 479
0 1156 5 1 1 483
0 1157 5 1 1 487
0 1158 6 1 2 1063 1064
0 1159 5 1 1 491
0 1160 6 1 2 492 892
0 1161 5 1 1 495
0 1162 6 1 2 1067 1068
0 1163 5 1 1 445
0 1164 1 2 1 446
0 1167 5 1 1 448
0 1168 1 2 1 449
0 1171 6 16 2 921 455
0 1188 6 16 2 922 456
0 1205 5 1 1 497
0 1206 6 1 2 498 938
0 1207 5 1 1 499
0 1208 6 1 2 500 942
0 1209 5 1 1 501
0 1210 6 1 2 502 946
0 1211 5 1 1 503
0 1212 6 1 2 504 950
0 1213 5 1 1 505
0 1214 6 1 2 506 954
0 1215 5 1 1 507
0 1216 6 1 2 508 958
0 1217 5 1 1 509
0 1218 5 1 1 477
0 1219 5 1 1 511
0 1220 5 1 1 513
0 1221 6 1 2 514 968
0 1222 5 1 1 481
0 1223 5 1 1 515
0 1224 6 1 2 516 972
0 1225 5 1 1 517
0 1226 6 1 2 518 976
0 1227 5 1 1 485
0 1228 5 1 1 519
0 1229 6 1 2 520 980
0 1230 5 1 1 489
0 1231 6 1 2 490 984
0 1232 6 2 2 1119 1120
0 1235 6 2 2 1121 1122
0 1238 5 1 1 521
0 1239 6 1 2 522 997
0 1240 5 1 1 493
0 1241 5 1 1 523
0 1242 6 1 2 524 1001
0 1243 6 2 2 1128 1129
0 1246 6 2 2 1130 1131
0 1249 6 2 2 1132 1133
0 1252 1 2 1 451
0 1255 1 2 1 452
0 1258 1 2 1 453
0 1261 1 2 1 454
0 1264 5 2 1 1150
0 1267 6 1 2 351 1159
0 1309 6 1 2 402 1205
0 1310 6 1 2 404 1207
0 1311 6 1 2 406 1209
0 1312 6 1 2 408 1211
0 1313 6 1 2 410 1213
0 1314 6 1 2 412 1215
0 1315 6 1 2 414 1220
0 1316 6 1 2 416 1223
0 1317 6 1 2 418 1225
0 1318 6 1 2 420 1228
0 1319 5 2 1 1158
0 1322 6 1 2 348 1230
0 1327 6 1 2 430 1238
0 1328 6 1 2 432 1241
0 1334 5 2 1 1162
0 1344 6 1 2 1267 1160
0 1345 6 1 2 610 894
0 1346 5 1 1 611
0 1348 5 1 1 615
0 1349 5 1 1 613
0 1350 5 1 1 621
0 1351 5 1 1 618
0 1352 6 2 2 1309 1206
0 1355 6 2 2 1310 1208
0 1358 6 2 2 1311 1210
0 1361 6 2 2 1312 1212
0 1364 6 2 2 1313 1214
0 1367 6 2 2 1314 1216
0 1370 6 2 2 1315 1221
0 1373 6 2 2 1316 1224
0 1376 6 2 2 1317 1226
0 1379 6 2 2 1318 1229
0 1383 6 2 2 1322 1231
0 1386 5 1 1 597
0 1387 6 1 2 599 990
0 1388 5 1 1 600
0 1389 6 1 2 604 993
0 1390 6 2 2 1327 1239
0 1393 6 2 2 1328 1242
0 1396 5 1 1 605
0 1397 6 1 2 606 1004
0 1398 5 1 1 607
0 1399 6 1 2 609 1007
0 1409 5 1 1 627
0 1412 6 1 2 369 1346
0 1413 5 1 1 630
0 1416 1 2 1 624
0 1419 1 2 1 626
0 1433 6 1 2 354 1386
0 1434 6 1 2 357 1388
0 1438 6 1 2 360 1396
0 1439 6 1 2 366 1398
0 1440 5 2 1 1344
0 1443 6 1 2 636 1148
0 1444 5 1 1 638
0 1445 6 1 2 633 1149
0 1446 5 1 1 635
0 1447 6 1 2 639 1151
0 1448 5 1 1 641
0 1451 6 1 2 642 1152
0 1452 5 1 1 644
0 1453 6 1 2 648 1153
0 1454 5 1 1 650
0 1455 6 1 2 645 1154
0 1456 5 1 1 647
0 1457 6 1 2 654 1156
0 1458 5 1 1 656
0 1459 6 1 2 660 1157
0 1460 5 1 1 662
0 1461 5 1 1 663
0 1462 6 1 2 669 1161
0 1463 5 1 1 671
0 1464 6 1 2 1345 1412
0 1468 5 1 1 651
0 1469 6 1 2 653 1222
0 1470 5 1 1 657
0 1471 6 1 2 659 1227
0 1472 6 2 2 1387 1433
0 1475 5 1 1 666
0 1476 6 1 2 668 1240
0 1478 6 2 2 1389 1434
0 1481 6 2 2 1399 1439
0 1484 6 2 2 1397 1438
0 1487 6 1 2 468 1444
0 1488 6 1 2 466 1446
0 1489 6 1 2 470 1448
0 1490 5 1 1 675
0 1491 5 1 1 672
0 1492 6 1 2 472 1452
0 1493 6 1 2 476 1454
0 1494 6 1 2 474 1456
0 1495 6 1 2 484 1458
0 1496 6 1 2 488 1460
0 1498 6 1 2 496 1463
0 1499 5 1 1 678
0 1500 6 1 2 482 1468
0 1501 6 1 2 486 1470
0 1504 6 1 2 494 1475
0 1510 5 2 1 1464
0 1513 6 1 2 1443 1487
0 1514 6 2 2 1445 1488
0 1517 6 2 2 1447 1489
0 1520 6 1 2 1451 1492
0 1521 6 1 2 1453 1493
0 1522 6 3 2 1455 1494
0 1526 6 1 2 1457 1495
0 1527 6 1 2 1459 1496
0 1528 5 1 1 681
0 1529 6 1 2 1462 1498
0 1530 5 1 1 684
0 1531 5 1 1 687
0 1532 5 1 1 690
0 1534 6 2 2 1471 1501
0 1537 6 2 2 1469 1500
0 1540 6 2 2 1476 1504
0 1546 5 2 1 1513
0 1554 5 2 1 1521
0 1557 5 3 1 1526
0 1561 5 2 1 1520
0 1567 6 1 2 692 1531
0 1568 6 1 2 689 1532
0 1569 5 1 1 693
0 1571 5 2 1 1527
0 1576 5 2 1 1529
0 1588 1 2 1 702
0 1591 5 1 1 707
0 1593 5 1 1 710
0 1594 6 1 2 713 1530
0 1595 5 1 1 714
0 1596 6 2 2 1567 1568
0 1600 1 2 1 699
0 1603 1 2 1 701
0 1606 1 2 1 704
0 1609 1 2 1 705
0 1612 1 2 1 696
0 1615 1 2 1 698
0 1620 1 2 1 722
0 1623 1 2 1 719
0 1635 5 1 1 729
0 1636 6 1 2 686 1595
0 1638 6 1 2 732 1569
0 1639 5 1 1 734
0 1640 1 2 1 726
0 1643 1 2 1 728
0 1647 1 2 1 716
0 1651 1 2 1 717
0 1658 1 2 1 720
0 1661 1 2 1 723
0 1664 1 2 1 725
0 1671 6 1 2 738 893
0 1672 5 1 1 740
0 1675 5 1 1 741
0 1677 5 1 1 744
0 1678 6 1 2 747 1217
0 1679 5 1 1 749
0 1680 6 1 2 750 1219
0 1681 5 1 1 752
0 1682 5 1 1 753
0 1683 5 1 1 755
0 1685 6 2 2 1594 1636
0 1688 6 1 2 695 1639
0 1697 1 2 1 735
0 1701 1 2 1 737
0 1706 6 1 2 363 1672
0 1707 5 1 1 763
0 1708 6 1 2 765 1675
0 1709 5 1 1 766
0 1710 6 1 2 767 1677
0 1711 5 1 1 768
0 1712 6 1 2 510 1679
0 1713 6 1 2 512 1681
0 1714 1 2 1 757
0 1717 1 2 1 758
0 1720 6 1 2 769 1593
0 1721 5 1 1 770
0 1723 6 2 2 1638 1688
0 1727 5 1 1 771
0 1728 5 1 1 761
0 1730 5 1 1 773
0 1731 1 2 1 759
0 1734 1 2 1 760
0 1740 6 1 2 775 1528
0 1741 5 1 1 776
0 1742 6 2 2 1671 1706
0 1746 6 1 2 743 1709
0 1747 6 1 2 746 1711
0 1748 6 2 2 1678 1712
0 1751 6 2 2 1680 1713
0 1759 6 1 2 711 1721
0 1761 5 1 1 777
0 1762 6 1 2 778 1727
0 1763 5 1 1 779
0 1764 6 1 2 780 1730
0 1768 5 1 1 783
0 1769 6 1 2 683 1741
0 1772 6 1 2 785 1413
0 1773 5 1 1 786
0 1774 6 2 2 1708 1746
0 1777 6 2 2 1710 1747
0 1783 5 1 1 787
0 1784 6 1 2 788 1682
0 1785 5 1 1 781
0 1786 5 1 1 789
0 1787 6 1 2 790 1683
0 1788 6 2 2 1720 1759
0 1791 6 1 2 772 1761
0 1792 6 1 2 774 1763
0 1795 6 1 2 795 1155
0 1796 5 1 1 796
0 1798 6 2 2 1740 1769
0 1801 6 1 2 632 1773
0 1802 6 2 2 791 181
0 1807 5 1 1 793
0 1808 6 1 2 794 1218
0 1809 6 1 2 754 1783
0 1810 6 1 2 756 1786
0 1812 6 2 2 1791 1762
0 1815 6 2 2 1792 1764
0 1818 1 2 1 792
0 1821 6 1 2 799 1490
0 1822 5 1 1 800
0 1823 6 1 2 797 1491
0 1824 5 1 1 798
0 1825 6 1 2 480 1796
0 1826 6 1 2 801 1409
0 1827 5 1 1 802
0 1830 6 2 2 1772 1801
0 1837 6 1 2 478 1807
0 1838 6 2 2 1809 1784
0 1841 6 2 2 1810 1787
0 1848 6 1 2 677 1822
0 1849 6 1 2 674 1824
0 1850 6 1 2 1795 1825
0 1852 6 1 2 629 1827
0 1855 6 1 2 809 1707
0 1856 5 1 1 810
0 1857 5 1 1 811
0 1858 6 2 2 803 182
0 1864 5 1 1 807
0 1865 6 1 2 808 1728
0 1866 1 2 1 804
0 1869 1 2 1 805
0 1872 1 2 1 806
0 1875 6 2 2 1808 1837
0 1878 6 1 2 1821 1848
0 1879 6 2 2 1823 1849
0 1882 6 1 2 817 1768
0 1883 5 1 1 818
0 1884 6 1 2 1826 1852
0 1885 6 1 2 764 1856
0 1889 6 2 2 813 183
0 1895 5 1 1 815
0 1896 6 1 2 816 1785
0 1897 6 1 2 762 1864
0 1898 5 2 1 1850
0 1902 1 2 1 814
0 1910 5 1 1 1878
0 1911 6 1 2 784 1883
0 1912 5 1 1 1884
0 1913 6 1 2 1855 1885
0 1915 5 1 1 821
0 1919 6 1 2 825 919
0 1920 5 1 1 826
0 1921 6 1 2 823 920
0 1922 5 1 1 824
0 1923 5 1 1 827
0 1924 6 1 2 782 1895
0 1927 1 2 1 819
0 1930 1 2 1 820
0 1933 6 2 2 1865 1897
0 1936 6 1 2 1882 1911
0 1937 5 1 1 833
0 1938 5 1 1 835
0 1941 6 1 2 396 1920
0 1942 6 1 2 394 1922
0 1944 1 2 1 829
0 1947 5 2 1 1913
0 1950 1 2 1 831
0 1953 1 2 1 832
0 1958 1 2 1 830
0 1961 6 2 2 1896 1924
0 1965 7 2 2 1910 601
0 1968 7 2 2 602 1912
0 1975 6 1 2 839 917
0 1976 5 1 1 840
0 1977 6 1 2 837 918
0 1978 5 1 1 838
0 1979 6 1 2 1919 1941
0 1980 6 2 2 1921 1942
0 1985 5 1 1 841
0 1987 5 2 1 1936
0 1999 5 1 1 843
0 2000 6 1 2 844 1937
0 2002 5 1 1 845
0 2003 6 1 2 846 1499
0 2004 6 1 2 849 1350
0 2005 5 1 1 850
0 2006 6 1 2 847 1351
0 2007 5 1 1 848
0 2008 6 1 2 392 1976
0 2009 6 1 2 390 1978
0 2012 5 1 1 1979
0 2013 5 1 1 851
0 2014 6 1 2 852 1923
0 2015 5 1 1 853
0 2016 6 1 2 854 1635
0 2018 5 1 1 855
0 2019 5 1 1 857
0 2020 6 1 2 834 1999
0 2021 5 1 1 861
0 2022 6 1 2 862 1591
0 2023 6 1 2 680 2002
0 2024 6 1 2 623 2005
0 2025 6 1 2 620 2007
0 2026 6 1 2 1975 2008
0 2027 6 2 2 1977 2009
0 2030 5 2 1 859
0 2033 1 2 1 860
0 2036 6 1 2 828 2013
0 2037 6 1 2 731 2015
0 2038 6 1 2 2020 2000
0 2039 6 1 2 708 2021
0 2040 6 1 2 2023 2003
0 2041 6 1 2 2004 2024
0 2042 6 2 2 2006 2025
0 2047 5 1 1 2026
0 2052 6 2 2 2036 2014
0 2055 6 2 2 2037 2016
0 2060 5 1 1 2038
0 2061 6 1 2 2039 2022
0 2062 6 2 2 2040 184
0 2067 5 1 1 2041
0 2068 5 2 1 863
0 2071 1 2 1 864
0 2076 5 1 1 871
0 2077 5 1 1 873
0 2078 6 2 2 2060 185
0 2081 6 2 2 2061 186
0 2086 5 2 1 869
0 2089 1 2 1 870
0 2104 7 14 2 865 877
0 2119 7 9 2 867 878
0 2129 7 13 2 866 879
0 2143 7 4 2 868 880
0 2148 1 2 1 875
0 2151 1 2 1 876
0 2196 1 2 1 881
0 2199 1 2 1 882
0 2202 1 2 1 883
0 2205 1 2 1 884
0 2214 6 1 2 983 915
0 2215 5 1 1 986
0 2216 6 1 2 979 916
0 2217 5 1 1 982
0 2222 6 1 2 996 1348
0 2223 5 1 1 999
0 2224 6 1 2 987 1349
0 2225 5 1 1 995
0 2226 6 1 2 1012 913
0 2227 5 1 1 1014
0 2228 6 1 2 1000 914
0 2229 5 1 1 1011
0 2230 6 1 2 387 2215
0 2231 6 1 2 384 2217
0 2232 6 1 2 617 2223
0 2233 6 1 2 614 2225
0 2234 6 1 2 381 2227
0 2235 6 1 2 378 2229
0 2236 6 1 2 2214 2230
0 2237 6 2 2 2216 2231
0 2240 6 1 2 2222 2232
0 2241 6 2 2 2224 2233
0 2244 6 1 2 2226 2234
0 2245 6 2 2 2228 2235
0 2250 5 1 1 2236
0 2253 5 1 1 2240
0 2256 5 1 1 2244
0 2257 5 2 1 1015
0 2260 1 2 1 1017
0 2263 5 2 1 1018
0 2266 7 2 2 525 1020
0 2269 5 2 1 1021
0 2272 7 2 2 527 1023
0 2279 6 2 8 2067 2012 2047 2250 447 2256 2253 450
0 2286 1 10 1 1033
0 2297 1 15 1 1035
0 2315 1 10 1 1039
0 2326 1 13 1 1041
0 2340 7 12 2 885 1024
0 2353 7 7 2 901 1026
0 2361 7 13 2 900 1027
0 2375 7 8 2 902 1029
0 2384 7 1 4 233 1042 203 203
0 2385 7 1 2 1163 1030
0 2386 7 14 2 526 1032
0 2426 7 1 2 1167 1036
0 2427 7 16 2 528 1038
0 2537 6 2 5 1045 1078 1124 904 529
0 2540 6 2 5 1047 1079 1101 948 530
0 2543 6 2 5 1048 1080 1102 932 531
0 2546 6 2 5 1050 1081 1113 905 532
0 2549 6 2 5 1059 1082 1143 933 573
0 2552 6 2 5 1060 1088 1125 971 575
0 2555 6 2 5 1061 1089 1144 949 576
0 2558 7 2 5 1051 1083 1126 906 533
0 2561 7 2 5 1052 1084 1103 952 557
0 2564 7 2 5 1053 1085 1104 934 558
0 2567 7 2 5 1056 1086 1114 908 560
0 2570 7 2 5 1062 1087 1145 936 578
0 2573 7 2 5 1065 1090 1127 974 579
0 2576 7 2 5 1066 1091 1146 953 581
0 2594 6 2 5 1057 1185 1134 956 561
0 2597 6 2 5 1069 1186 1135 937 563
0 2600 6 2 5 1070 1187 1147 909 564
0 2603 6 2 5 1071 1189 1105 975 566
0 2606 6 2 5 1072 1190 1115 957 582
0 2611 6 2 5 1170 1092 1136 960 584
0 2614 6 2 5 1172 1093 1137 940 585
0 2617 6 2 5 1173 1094 1165 911 587
0 2620 6 2 5 1174 1095 1116 961 588
0 2627 6 1 5 1073 1191 1106 912 457
0 2628 6 1 5 1175 1096 1107 924 458
0 2629 6 1 5 1176 1192 1138 925 459
0 2630 6 1 5 1177 1193 1108 963 460
0 2631 6 1 5 1178 1194 1109 941 461
0 2632 6 1 5 1179 1195 1117 927 462
0 2633 6 1 5 1180 2426 1110 928 463
0 2634 6 1 5 2385 1196 1111 929 464
0 2639 7 2 5 1058 1197 1139 964 567
0 2642 7 2 5 1074 1198 1140 944 569
0 2645 7 2 5 1075 1199 1166 930 570
0 2648 7 2 5 1076 1200 1112 978 572
0 2651 7 2 5 1077 1201 1118 966 590
0 2655 7 2 5 1181 1097 1141 967 591
0 2658 7 2 5 1182 1098 1142 945 593
0 2661 7 2 5 1183 1099 1169 931 594
0 2664 7 2 5 1184 1100 1123 970 596
0 2669 6 1 2 1254 534
0 2670 5 1 1 1256
0 2671 6 1 2 1257 535
0 2672 5 1 1 1259
0 2673 6 1 2 1260 536
0 2674 5 1 1 1262
0 2675 6 1 2 1263 537
0 2676 5 1 1 1265
0 2682 6 1 2 1266 543
0 2683 5 1 1 1268
0 2688 6 1 2 1269 548
0 2689 5 1 1 1270
0 2690 6 1 2 1271 549
0 2691 5 1 1 1272
0 2710 7 1 8 2627 2628 2629 2630 2631 2632 2633 2634
0 2720 6 1 2 237 2670
0 2721 6 1 2 240 2672
0 2722 6 1 2 242 2674
0 2723 6 1 2 245 2676
0 2724 6 1 2 1291 538
0 2725 5 1 1 1292
0 2726 6 1 2 1293 539
0 2727 5 1 1 1294
0 2728 6 1 2 1295 540
0 2729 5 1 1 1296
0 2730 6 1 2 1297 541
0 2731 5 1 1 1298
0 2732 6 1 2 1299 542
0 2733 5 1 1 1300
0 2734 6 1 2 265 2683
0 2735 6 1 2 1301 544
0 2736 5 1 1 1302
0 2737 6 1 2 1303 545
0 2738 5 1 1 1304
0 2739 6 1 2 1305 546
0 2740 5 1 1 1306
0 2741 6 1 2 1307 547
0 2742 5 1 1 1308
0 2743 6 1 2 282 2689
0 2744 6 1 2 285 2691
0 2745 6 1 8 1202 1204 1234 1237 1273 1275 1277 1279
0 2746 6 1 8 1281 1245 1283 1285 1287 1289 1248 1251
0 2747 7 2 8 1203 1233 1236 1244 1274 1276 1278 1280
0 2750 7 2 8 1282 1247 1284 1286 1288 1290 1250 1253
3 2753 6 0 2 2669 2720
3 2754 6 0 2 2671 2721
3 2755 6 0 2 2673 2722
3 2756 6 0 2 2675 2723
0 2757 6 1 2 248 2725
0 2758 6 1 2 250 2727
0 2759 6 1 2 255 2729
0 2760 6 1 2 259 2731
0 2761 6 1 2 262 2733
3 2762 6 0 2 2682 2734
0 2763 6 1 2 268 2736
0 2764 6 1 2 271 2738
0 2765 6 1 2 274 2740
0 2766 6 1 2 279 2742
3 2767 6 0 2 2688 2743
3 2768 6 0 2 2690 2744
0 2773 7 2 2 2745 275
0 2776 7 2 2 2746 276
3 2779 6 0 2 2724 2757
3 2780 6 0 2 2726 2758
3 2781 6 0 2 2728 2759
3 2782 6 0 2 2730 2760
3 2783 6 0 2 2732 2761
3 2784 6 0 2 2735 2763
3 2785 6 0 2 2737 2764
3 2786 6 0 2 2739 2765
3 2787 6 0 2 2741 2766
0 2788 7 1 3 1320 1323 2710
0 2789 6 6 2 1321 1324
0 2800 7 1 4 234 1044 103 2788
0 2807 6 1 2 1325 2018
0 2808 5 1 1 1326
0 2809 6 1 2 1329 2019
0 2810 5 1 1 1330
3 2811 4 0 2 2384 2800
0 2812 7 2 3 897 175 1331
0 2815 7 2 3 78 176 1332
0 2818 7 2 3 84 177 1333
0 2821 7 2 3 87 178 1335
0 2824 7 2 3 898 179 1336
0 2827 6 1 2 856 2808
0 2828 6 1 2 858 2810
0 2829 7 2 3 81 180 1337
0 2843 6 2 2 2807 2827
0 2846 6 2 2 2809 2828
0 2850 6 1 2 1338 2076
0 2851 6 1 2 1340 2077
0 2852 6 1 2 1342 1915
0 2853 6 1 2 1347 1857
0 2854 6 1 2 1354 1938
0 2857 5 1 1 1339
0 2858 5 1 1 1341
0 2859 5 1 1 1343
0 2860 5 1 1 1353
0 2861 5 1 1 1356
0 2862 5 1 1 1357
0 2863 6 1 2 1359 1985
0 2866 6 1 2 872 2857
0 2867 6 1 2 874 2858
0 2868 6 1 2 822 2859
0 2869 6 1 2 812 2860
0 2870 6 1 2 836 2861
0 2871 6 1 2 1360 886
0 2872 5 1 1 1362
0 2873 6 1 2 1363 887
0 2874 5 1 1 1365
0 2875 6 1 2 842 2862
0 2876 6 1 2 2866 2850
0 2877 6 1 2 2867 2851
0 2878 6 1 2 2868 2852
0 2879 6 1 2 2869 2853
0 2880 6 1 2 2870 2854
0 2881 6 1 2 398 2872
0 2882 6 1 2 400 2874
0 2883 6 2 2 2875 2863
3 2886 7 0 2 2876 550
3 2887 7 0 2 551 2877
3 2888 7 0 2 553 2878
3 2889 7 0 2 2879 554
3 2890 7 0 2 555 2880
3 2891 6 0 2 2871 2881
3 2892 6 0 2 2873 2882
0 2895 6 1 2 1366 1461
0 2896 5 1 1 1368
0 2897 6 1 2 665 2896
0 2898 6 1 2 2895 2897
3 2899 7 0 2 2898 552
2 2 1 1
2 3 1 1
2 5 1 4
2 6 1 4
2 8 1 7
2 9 1 7
2 11 1 10
2 12 1 10
2 14 1 13
2 15 1 13
2 17 1 16
2 18 1 16
2 20 1 19
2 21 1 19
2 23 1 22
2 24 1 22
2 26 1 25
2 27 1 25
2 29 1 28
2 30 1 28
2 32 1 31
2 33 1 31
2 35 1 34
2 36 1 34
2 38 1 37
2 39 1 37
2 41 1 40
2 42 1 40
2 44 1 43
2 45 1 43
2 47 1 46
2 48 1 46
2 50 1 49
2 51 1 49
2 52 1 49
2 54 1 53
2 55 1 53
2 57 1 56
2 58 1 56
2 59 1 56
2 61 1 60
2 62 1 60
2 64 1 63
2 65 1 63
2 67 1 66
2 68 1 66
2 70 1 69
2 71 1 69
2 73 1 72
2 74 1 72
2 75 1 72
2 77 1 76
2 78 1 76
2 80 1 79
2 81 1 79
2 83 1 82
2 84 1 82
2 86 1 85
2 87 1 85
2 89 1 88
2 90 1 88
2 92 1 91
2 93 1 91
2 95 1 94
2 96 1 94
2 97 1 94
2 98 1 94
2 100 1 99
2 101 1 99
2 102 1 99
2 103 1 99
2 105 1 104
2 106 1 104
2 107 1 104
2 108 1 104
2 109 1 104
2 110 1 104
2 111 1 104
2 112 1 190
2 113 1 190
2 114 1 190
2 115 1 194
2 116 1 194
2 117 1 197
2 118 1 197
2 119 1 197
2 120 1 201
2 121 1 201
2 122 1 201
2 123 1 201
2 124 1 206
2 125 1 206
2 126 1 209
2 127 1 209
2 128 1 212
2 129 1 212
2 130 1 212
2 131 1 216
2 132 1 216
2 133 1 216
2 134 1 220
2 135 1 220
2 136 1 220
2 137 1 220
2 138 1 225
2 139 1 225
2 140 1 225
2 141 1 229
2 142 1 229
2 143 1 232
2 144 1 232
2 145 1 235
2 146 1 235
2 147 1 235
2 148 1 239
2 149 1 239
2 150 1 239
2 151 1 243
2 152 1 243
2 153 1 243
2 154 1 247
2 155 1 247
2 156 1 247
2 157 1 253
2 158 1 253
2 159 1 257
2 160 1 257
2 161 1 260
2 162 1 260
2 163 1 263
2 164 1 263
2 165 1 266
2 166 1 266
2 167 1 269
2 168 1 269
2 169 1 272
2 170 1 272
2 171 1 277
2 172 1 277
2 173 1 280
2 174 1 280
2 175 1 283
2 176 1 283
2 177 1 283
2 178 1 283
2 179 1 283
2 180 1 283
2 181 1 290
2 182 1 290
2 183 1 290
2 184 1 290
2 185 1 290
2 186 1 290
2 187 1 297
2 188 1 297
2 189 1 300
2 191 1 300
2 192 1 303
2 193 1 303
2 195 1 306
2 196 1 306
2 198 1 306
2 199 1 306
2 200 1 306
2 202 1 306
2 203 1 313
2 204 1 313
2 205 1 316
2 207 1 316
2 208 1 319
2 210 1 319
2 211 1 319
2 213 1 319
2 214 1 319
2 215 1 319
2 217 1 326
2 218 1 326
2 219 1 326
2 221 1 326
2 222 1 331
2 223 1 331
2 224 1 331
2 226 1 331
2 227 1 331
2 228 1 331
2 230 1 338
2 231 1 338
2 233 1 338
2 234 1 338
2 236 1 343
2 237 1 343
2 238 1 346
2 240 1 346
2 241 1 349
2 242 1 349
2 244 1 352
2 245 1 352
2 246 1 355
2 248 1 355
2 249 1 358
2 250 1 358
2 254 1 361
2 255 1 361
2 258 1 364
2 259 1 364
2 261 1 367
2 262 1 367
2 264 1 370
2 265 1 370
2 267 1 373
2 268 1 373
2 270 1 376
2 271 1 376
2 273 1 379
2 274 1 379
2 278 1 382
2 279 1 382
2 281 1 385
2 282 1 385
2 284 1 388
2 285 1 388
2 286 1 556
2 287 1 556
2 288 1 559
2 289 1 559
2 291 1 562
2 292 1 562
2 293 1 565
2 294 1 565
2 295 1 568
2 296 1 568
2 298 1 571
2 299 1 571
2 301 1 574
2 302 1 574
2 304 1 577
2 305 1 577
2 307 1 580
2 308 1 580
2 309 1 583
2 310 1 583
2 311 1 586
2 312 1 586
2 314 1 589
2 315 1 589
2 317 1 592
2 318 1 592
2 320 1 595
2 321 1 595
2 322 1 598
2 323 1 598
2 324 1 603
2 325 1 603
2 327 1 603
2 328 1 603
2 329 1 608
2 330 1 608
2 332 1 608
2 333 1 612
2 334 1 612
2 335 1 612
2 336 1 616
2 337 1 616
2 339 1 619
2 340 1 619
2 341 1 622
2 342 1 622
2 344 1 625
2 345 1 625
2 347 1 628
2 348 1 628
2 350 1 631
2 351 1 631
2 353 1 634
2 354 1 634
2 356 1 637
2 357 1 637
2 359 1 640
2 360 1 640
2 362 1 643
2 363 1 643
2 365 1 646
2 366 1 646
2 368 1 649
2 369 1 649
2 371 1 652
2 372 1 652
2 374 1 655
2 375 1 655
2 377 1 658
2 378 1 658
2 380 1 661
2 381 1 661
2 383 1 664
2 384 1 664
2 386 1 667
2 387 1 667
2 389 1 670
2 390 1 670
2 391 1 673
2 392 1 673
2 393 1 676
2 394 1 676
2 395 1 679
2 396 1 679
2 397 1 682
2 398 1 682
2 399 1 685
2 400 1 685
2 401 1 688
2 402 1 688
2 403 1 691
2 404 1 691
2 405 1 694
2 406 1 694
2 407 1 697
2 408 1 697
2 409 1 700
2 410 1 700
2 411 1 703
2 412 1 703
2 413 1 706
2 414 1 706
2 415 1 709
2 416 1 709
2 417 1 712
2 418 1 712
2 419 1 715
2 420 1 715
2 421 1 718
2 422 1 718
2 423 1 721
2 424 1 721
2 425 1 724
2 426 1 724
2 427 1 727
2 428 1 727
2 429 1 730
2 430 1 730
2 431 1 733
2 432 1 733
2 433 1 736
2 434 1 736
2 435 1 739
2 436 1 739
2 437 1 742
2 438 1 742
2 439 1 745
2 440 1 745
2 441 1 748
2 442 1 748
2 443 1 751
2 444 1 751
2 445 1 899
2 446 1 899
2 447 1 899
2 448 1 903
2 449 1 903
2 450 1 903
2 451 1 907
2 452 1 907
2 453 1 910
2 454 1 910
2 455 1 923
2 456 1 923
2 457 1 926
2 458 1 926
2 459 1 926
2 460 1 926
2 461 1 926
2 462 1 926
2 463 1 926
2 464 1 926
2 465 1 935
2 466 1 935
2 467 1 939
2 468 1 939
2 469 1 943
2 470 1 943
2 471 1 947
2 472 1 947
2 473 1 951
2 474 1 951
2 475 1 955
2 476 1 955
2 477 1 959
2 478 1 959
2 479 1 962
2 480 1 962
2 481 1 965
2 482 1 965
2 483 1 969
2 484 1 969
2 485 1 973
2 486 1 973
2 487 1 977
2 488 1 977
2 489 1 981
2 490 1 981
2 491 1 985
2 492 1 985
2 493 1 994
2 494 1 994
2 495 1 998
2 496 1 998
2 497 1 1010
2 498 1 1010
2 499 1 1013
2 500 1 1013
2 501 1 1016
2 502 1 1016
2 503 1 1019
2 504 1 1019
2 505 1 1022
2 506 1 1022
2 507 1 1025
2 508 1 1025
2 509 1 1028
2 510 1 1028
2 511 1 1031
2 512 1 1031
2 513 1 1034
2 514 1 1034
2 515 1 1037
2 516 1 1037
2 517 1 1040
2 518 1 1040
2 519 1 1043
2 520 1 1043
2 521 1 1046
2 522 1 1046
2 523 1 1049
2 524 1 1049
2 525 1 1164
2 526 1 1164
2 527 1 1168
2 528 1 1168
2 529 1 1171
2 530 1 1171
2 531 1 1171
2 532 1 1171
2 533 1 1171
2 557 1 1171
2 558 1 1171
2 560 1 1171
2 561 1 1171
2 563 1 1171
2 564 1 1171
2 566 1 1171
2 567 1 1171
2 569 1 1171
2 570 1 1171
2 572 1 1171
2 573 1 1188
2 575 1 1188
2 576 1 1188
2 578 1 1188
2 579 1 1188
2 581 1 1188
2 582 1 1188
2 584 1 1188
2 585 1 1188
2 587 1 1188
2 588 1 1188
2 590 1 1188
2 591 1 1188
2 593 1 1188
2 594 1 1188
2 596 1 1188
2 597 1 1232
2 599 1 1232
2 600 1 1235
2 604 1 1235
2 605 1 1243
2 606 1 1243
2 607 1 1246
2 609 1 1246
2 610 1 1249
2 611 1 1249
2 613 1 1252
2 614 1 1252
2 615 1 1255
2 617 1 1255
2 618 1 1258
2 620 1 1258
2 621 1 1261
2 623 1 1261
2 624 1 1264
2 626 1 1264
2 627 1 1319
2 629 1 1319
2 630 1 1334
2 632 1 1334
2 633 1 1352
2 635 1 1352
2 636 1 1355
2 638 1 1355
2 639 1 1358
2 641 1 1358
2 642 1 1361
2 644 1 1361
2 645 1 1364
2 647 1 1364
2 648 1 1367
2 650 1 1367
2 651 1 1370
2 653 1 1370
2 654 1 1373
2 656 1 1373
2 657 1 1376
2 659 1 1376
2 660 1 1379
2 662 1 1379
2 663 1 1383
2 665 1 1383
2 666 1 1390
2 668 1 1390
2 669 1 1393
2 671 1 1393
2 672 1 1416
2 674 1 1416
2 675 1 1419
2 677 1 1419
2 678 1 1440
2 680 1 1440
2 681 1 1472
2 683 1 1472
2 684 1 1478
2 686 1 1478
2 687 1 1481
2 689 1 1481
2 690 1 1484
2 692 1 1484
2 693 1 1510
2 695 1 1510
2 696 1 1514
2 698 1 1514
2 699 1 1517
2 701 1 1517
2 702 1 1522
2 704 1 1522
2 705 1 1522
2 707 1 1534
2 708 1 1534
2 710 1 1537
2 711 1 1537
2 713 1 1540
2 714 1 1540
2 716 1 1546
2 717 1 1546
2 719 1 1554
2 720 1 1554
2 722 1 1557
2 723 1 1557
2 725 1 1557
2 726 1 1561
2 728 1 1561
2 729 1 1571
2 731 1 1571
2 732 1 1576
2 734 1 1576
2 735 1 1588
2 737 1 1588
2 738 1 1596
2 740 1 1596
2 741 1 1600
2 743 1 1600
2 744 1 1603
2 746 1 1603
2 747 1 1606
2 749 1 1606
2 750 1 1609
2 752 1 1609
2 753 1 1612
2 754 1 1612
2 755 1 1615
2 756 1 1615
2 757 1 1620
2 758 1 1620
2 759 1 1623
2 760 1 1623
2 761 1 1640
2 762 1 1640
2 763 1 1643
2 764 1 1643
2 765 1 1647
2 766 1 1647
2 767 1 1651
2 768 1 1651
2 769 1 1658
2 770 1 1658
2 771 1 1661
2 772 1 1661
2 773 1 1664
2 774 1 1664
2 775 1 1685
2 776 1 1685
2 777 1 1697
2 778 1 1697
2 779 1 1701
2 780 1 1701
2 781 1 1714
2 782 1 1714
2 783 1 1717
2 784 1 1717
2 785 1 1723
2 786 1 1723
2 787 1 1731
2 788 1 1731
2 789 1 1734
2 790 1 1734
2 791 1 1742
2 792 1 1742
2 793 1 1748
2 794 1 1748
2 795 1 1751
2 796 1 1751
2 797 1 1774
2 798 1 1774
2 799 1 1777
2 800 1 1777
2 801 1 1788
2 802 1 1788
2 803 1 1798
2 804 1 1798
2 805 1 1802
2 806 1 1802
2 807 1 1812
2 808 1 1812
2 809 1 1815
2 810 1 1815
2 811 1 1818
2 812 1 1818
2 813 1 1830
2 814 1 1830
2 815 1 1838
2 816 1 1838
2 817 1 1841
2 818 1 1841
2 819 1 1858
2 820 1 1858
2 821 1 1866
2 822 1 1866
2 823 1 1869
2 824 1 1869
2 825 1 1872
2 826 1 1872
2 827 1 1875
2 828 1 1875
2 829 1 1879
2 830 1 1879
2 831 1 1889
2 832 1 1889
2 833 1 1898
2 834 1 1898
2 835 1 1902
2 836 1 1902
2 837 1 1927
2 838 1 1927
2 839 1 1930
2 840 1 1930
2 841 1 1933
2 842 1 1933
2 843 1 1944
2 844 1 1944
2 845 1 1947
2 846 1 1947
2 847 1 1950
2 848 1 1950
2 849 1 1953
2 850 1 1953
2 851 1 1958
2 852 1 1958
2 853 1 1961
2 854 1 1961
2 855 1 1965
2 856 1 1965
2 857 1 1968
2 858 1 1968
2 859 1 1980
2 860 1 1980
2 861 1 1987
2 862 1 1987
2 863 1 2027
2 864 1 2027
2 865 1 2030
2 866 1 2030
2 867 1 2033
2 868 1 2033
2 869 1 2042
2 870 1 2042
2 871 1 2052
2 872 1 2052
2 873 1 2055
2 874 1 2055
2 875 1 2062
2 876 1 2062
2 877 1 2068
2 878 1 2068
2 879 1 2071
2 880 1 2071
2 881 1 2078
2 882 1 2078
2 883 1 2081
2 884 1 2081
2 885 1 2086
2 900 1 2086
2 901 1 2089
2 902 1 2089
2 904 1 2104
2 905 1 2104
2 906 1 2104
2 908 1 2104
2 909 1 2104
2 911 1 2104
2 912 1 2104
2 924 1 2104
2 925 1 2104
2 927 1 2104
2 928 1 2104
2 929 1 2104
2 930 1 2104
2 931 1 2104
2 932 1 2119
2 933 1 2119
2 934 1 2119
2 936 1 2119
2 937 1 2119
2 940 1 2119
2 941 1 2119
2 944 1 2119
2 945 1 2119
2 948 1 2129
2 949 1 2129
2 952 1 2129
2 953 1 2129
2 956 1 2129
2 957 1 2129
2 960 1 2129
2 961 1 2129
2 963 1 2129
2 964 1 2129
2 966 1 2129
2 967 1 2129
2 970 1 2129
2 971 1 2143
2 974 1 2143
2 975 1 2143
2 978 1 2143
2 979 1 2148
2 982 1 2148
2 983 1 2151
2 986 1 2151
2 987 1 2196
2 995 1 2196
2 996 1 2199
2 999 1 2199
2 1000 1 2202
2 1011 1 2202
2 1012 1 2205
2 1014 1 2205
2 1015 1 2237
2 1017 1 2237
2 1018 1 2241
2 1020 1 2241
2 1021 1 2245
2 1023 1 2245
2 1024 1 2257
2 1026 1 2257
2 1027 1 2260
2 1029 1 2260
2 1030 1 2263
2 1032 1 2263
2 1033 1 2266
2 1035 1 2266
2 1036 1 2269
2 1038 1 2269
2 1039 1 2272
2 1041 1 2272
2 1042 1 2279
2 1044 1 2279
2 1045 1 2286
2 1047 1 2286
2 1048 1 2286
2 1050 1 2286
2 1051 1 2286
2 1052 1 2286
2 1053 1 2286
2 1056 1 2286
2 1057 1 2286
2 1058 1 2286
2 1059 1 2297
2 1060 1 2297
2 1061 1 2297
2 1062 1 2297
2 1065 1 2297
2 1066 1 2297
2 1069 1 2297
2 1070 1 2297
2 1071 1 2297
2 1072 1 2297
2 1073 1 2297
2 1074 1 2297
2 1075 1 2297
2 1076 1 2297
2 1077 1 2297
2 1078 1 2315
2 1079 1 2315
2 1080 1 2315
2 1081 1 2315
2 1082 1 2315
2 1083 1 2315
2 1084 1 2315
2 1085 1 2315
2 1086 1 2315
2 1087 1 2315
2 1088 1 2326
2 1089 1 2326
2 1090 1 2326
2 1091 1 2326
2 1092 1 2326
2 1093 1 2326
2 1094 1 2326
2 1095 1 2326
2 1096 1 2326
2 1097 1 2326
2 1098 1 2326
2 1099 1 2326
2 1100 1 2326
2 1101 1 2340
2 1102 1 2340
2 1103 1 2340
2 1104 1 2340
2 1105 1 2340
2 1106 1 2340
2 1107 1 2340
2 1108 1 2340
2 1109 1 2340
2 1110 1 2340
2 1111 1 2340
2 1112 1 2340
2 1113 1 2353
2 1114 1 2353
2 1115 1 2353
2 1116 1 2353
2 1117 1 2353
2 1118 1 2353
2 1123 1 2353
2 1124 1 2361
2 1125 1 2361
2 1126 1 2361
2 1127 1 2361
2 1134 1 2361
2 1135 1 2361
2 1136 1 2361
2 1137 1 2361
2 1138 1 2361
2 1139 1 2361
2 1140 1 2361
2 1141 1 2361
2 1142 1 2361
2 1143 1 2375
2 1144 1 2375
2 1145 1 2375
2 1146 1 2375
2 1147 1 2375
2 1165 1 2375
2 1166 1 2375
2 1169 1 2375
2 1170 1 2386
2 1172 1 2386
2 1173 1 2386
2 1174 1 2386
2 1175 1 2386
2 1176 1 2386
2 1177 1 2386
2 1178 1 2386
2 1179 1 2386
2 1180 1 2386
2 1181 1 2386
2 1182 1 2386
2 1183 1 2386
2 1184 1 2386
2 1185 1 2427
2 1186 1 2427
2 1187 1 2427
2 1189 1 2427
2 1190 1 2427
2 1191 1 2427
2 1192 1 2427
2 1193 1 2427
2 1194 1 2427
2 1195 1 2427
2 1196 1 2427
2 1197 1 2427
2 1198 1 2427
2 1199 1 2427
2 1200 1 2427
2 1201 1 2427
2 1202 1 2537
2 1203 1 2537
2 1204 1 2540
2 1233 1 2540
2 1234 1 2543
2 1236 1 2543
2 1237 1 2546
2 1244 1 2546
2 1245 1 2549
2 1247 1 2549
2 1248 1 2552
2 1250 1 2552
2 1251 1 2555
2 1253 1 2555
2 1254 1 2558
2 1256 1 2558
2 1257 1 2561
2 1259 1 2561
2 1260 1 2564
2 1262 1 2564
2 1263 1 2567
2 1265 1 2567
2 1266 1 2570
2 1268 1 2570
2 1269 1 2573
2 1270 1 2573
2 1271 1 2576
2 1272 1 2576
2 1273 1 2594
2 1274 1 2594
2 1275 1 2597
2 1276 1 2597
2 1277 1 2600
2 1278 1 2600
2 1279 1 2603
2 1280 1 2603
2 1281 1 2606
2 1282 1 2606
2 1283 1 2611
2 1284 1 2611
2 1285 1 2614
2 1286 1 2614
2 1287 1 2617
2 1288 1 2617
2 1289 1 2620
2 1290 1 2620
2 1291 1 2639
2 1292 1 2639
2 1293 1 2642
2 1294 1 2642
2 1295 1 2645
2 1296 1 2645
2 1297 1 2648
2 1298 1 2648
2 1299 1 2651
2 1300 1 2651
2 1301 1 2655
2 1302 1 2655
2 1303 1 2658
2 1304 1 2658
2 1305 1 2661
2 1306 1 2661
2 1307 1 2664
2 1308 1 2664
2 1320 1 2747
2 1321 1 2747
2 1323 1 2750
2 1324 1 2750
2 1325 1 2773
2 1326 1 2773
2 1329 1 2776
2 1330 1 2776
2 1331 1 2789
2 1332 1 2789
2 1333 1 2789
2 1335 1 2789
2 1336 1 2789
2 1337 1 2789
2 1338 1 2812
2 1339 1 2812
2 1340 1 2815
2 1341 1 2815
2 1342 1 2818
2 1343 1 2818
2 1347 1 2821
2 1353 1 2821
2 1354 1 2824
2 1356 1 2824
2 1357 1 2829
2 1359 1 2829
2 1360 1 2843
2 1362 1 2843
2 1363 1 2846
2 1365 1 2846
2 1366 1 2883
2 1368 1 2883
