1 1 0 6 0
1 8 0 6 0
1 15 0 6 0
1 22 0 6 0
1 29 0 6 0
1 36 0 6 0
1 43 0 6 0
1 50 0 6 0
1 57 0 6 0
1 64 0 6 0
1 71 0 6 0
1 78 0 6 0
1 85 0 6 0
1 92 0 6 0
1 99 0 6 0
1 106 0 6 0
1 113 0 6 0
1 120 0 6 0
1 127 0 6 0
1 134 0 6 0
1 141 0 6 0
1 148 0 6 0
1 155 0 6 0
1 162 0 6 0
1 169 0 6 0
1 176 0 6 0
1 183 0 6 0
1 190 0 6 0
1 197 0 6 0
1 204 0 6 0
1 211 0 6 0
1 218 0 6 0
1 225 0 1 0
1 226 0 1 0
1 227 0 1 0
1 228 0 1 0
1 229 0 1 0
1 230 0 1 0
1 231 0 1 0
1 232 0 1 0
1 233 0 8 0
0 242 7 2 2 225 234
0 245 7 2 2 226 235
0 248 7 2 2 227 236
0 251 7 2 2 228 237
0 254 7 2 2 229 238
0 257 7 2 2 230 239
0 260 7 2 2 231 240
0 263 7 2 2 232 241
0 266 6 2 2 2 9
0 269 6 2 2 16 23
0 272 6 2 2 30 37
0 275 6 2 2 44 51
0 278 6 2 2 58 65
0 281 6 2 2 72 79
0 284 6 2 2 86 93
0 287 6 2 2 100 107
0 290 6 2 2 114 121
0 293 6 2 2 128 135
0 296 6 2 2 142 149
0 299 6 2 2 156 163
0 302 6 2 2 170 177
0 305 6 2 2 184 191
0 308 6 2 2 198 205
0 311 6 2 2 212 219
0 314 6 2 2 3 31
0 317 6 2 2 59 87
0 320 6 2 2 10 38
0 323 6 2 2 66 94
0 326 6 2 2 17 45
0 329 6 2 2 73 101
0 332 6 2 2 24 52
0 335 6 2 2 80 108
0 338 6 2 2 115 143
0 341 6 2 2 171 199
0 344 6 2 2 122 150
0 347 6 2 2 178 206
0 350 6 2 2 129 157
0 353 6 2 2 185 213
0 356 6 2 2 136 164
0 359 6 2 2 192 220
0 362 6 1 2 4 267
0 363 6 1 2 11 268
0 364 6 1 2 18 270
0 365 6 1 2 25 271
0 366 6 1 2 32 273
0 367 6 1 2 39 274
0 368 6 1 2 46 276
0 369 6 1 2 53 277
0 370 6 1 2 60 279
0 371 6 1 2 67 280
0 372 6 1 2 74 282
0 373 6 1 2 81 283
0 374 6 1 2 88 285
0 375 6 1 2 95 286
0 376 6 1 2 102 288
0 377 6 1 2 109 289
0 378 6 1 2 116 291
0 379 6 1 2 123 292
0 380 6 1 2 130 294
0 381 6 1 2 137 295
0 382 6 1 2 144 297
0 383 6 1 2 151 298
0 384 6 1 2 158 300
0 385 6 1 2 165 301
0 386 6 1 2 172 303
0 387 6 1 2 179 304
0 388 6 1 2 186 306
0 389 6 1 2 193 307
0 390 6 1 2 200 309
0 391 6 1 2 207 310
0 392 6 1 2 214 312
0 393 6 1 2 221 313
0 394 6 1 2 5 315
0 395 6 1 2 33 316
0 396 6 1 2 61 318
0 397 6 1 2 89 319
0 398 6 1 2 12 321
0 399 6 1 2 40 322
0 400 6 1 2 68 324
0 401 6 1 2 96 325
0 402 6 1 2 19 327
0 403 6 1 2 47 328
0 404 6 1 2 75 330
0 405 6 1 2 103 331
0 406 6 1 2 26 333
0 407 6 1 2 54 334
0 408 6 1 2 82 336
0 409 6 1 2 110 337
0 410 6 1 2 117 339
0 411 6 1 2 145 340
0 412 6 1 2 173 342
0 413 6 1 2 201 343
0 414 6 1 2 124 345
0 415 6 1 2 152 346
0 416 6 1 2 180 348
0 417 6 1 2 208 349
0 418 6 1 2 131 351
0 419 6 1 2 159 352
0 420 6 1 2 187 354
0 421 6 1 2 215 355
0 422 6 1 2 138 357
0 423 6 1 2 166 358
0 424 6 1 2 194 360
0 425 6 1 2 222 361
0 426 6 2 2 362 363
0 429 6 2 2 364 365
0 432 6 2 2 366 367
0 435 6 2 2 368 369
0 438 6 2 2 370 371
0 441 6 2 2 372 373
0 444 6 2 2 374 375
0 447 6 2 2 376 377
0 450 6 2 2 378 379
0 453 6 2 2 380 381
0 456 6 2 2 382 383
0 459 6 2 2 384 385
0 462 6 2 2 386 387
0 465 6 2 2 388 389
0 468 6 2 2 390 391
0 471 6 2 2 392 393
0 474 6 2 2 394 395
0 477 6 2 2 396 397
0 480 6 2 2 398 399
0 483 6 2 2 400 401
0 486 6 2 2 402 403
0 489 6 2 2 404 405
0 492 6 2 2 406 407
0 495 6 2 2 408 409
0 498 6 2 2 410 411
0 501 6 2 2 412 413
0 504 6 2 2 414 415
0 507 6 2 2 416 417
0 510 6 2 2 418 419
0 513 6 2 2 420 421
0 516 6 2 2 422 423
0 519 6 2 2 424 425
0 522 6 2 2 427 430
0 525 6 2 2 433 436
0 528 6 2 2 439 442
0 531 6 2 2 445 448
0 534 6 2 2 451 454
0 537 6 2 2 457 460
0 540 6 2 2 463 466
0 543 6 2 2 469 472
0 546 6 2 2 475 478
0 549 6 2 2 481 484
0 552 6 2 2 487 490
0 555 6 2 2 493 496
0 558 6 2 2 499 502
0 561 6 2 2 505 508
0 564 6 2 2 511 514
0 567 6 2 2 517 520
0 570 6 1 2 428 523
0 571 6 1 2 431 524
0 572 6 1 2 434 526
0 573 6 1 2 437 527
0 574 6 1 2 440 529
0 575 6 1 2 443 530
0 576 6 1 2 446 532
0 577 6 1 2 449 533
0 578 6 1 2 452 535
0 579 6 1 2 455 536
0 580 6 1 2 458 538
0 581 6 1 2 461 539
0 582 6 1 2 464 541
0 583 6 1 2 467 542
0 584 6 1 2 470 544
0 585 6 1 2 473 545
0 586 6 1 2 476 547
0 587 6 1 2 479 548
0 588 6 1 2 482 550
0 589 6 1 2 485 551
0 590 6 1 2 488 553
0 591 6 1 2 491 554
0 592 6 1 2 494 556
0 593 6 1 2 497 557
0 594 6 1 2 500 559
0 595 6 1 2 503 560
0 596 6 1 2 506 562
0 597 6 1 2 509 563
0 598 6 1 2 512 565
0 599 6 1 2 515 566
0 600 6 1 2 518 568
0 601 6 1 2 521 569
0 602 6 4 2 570 571
0 607 6 4 2 572 573
0 612 6 4 2 574 575
0 617 6 4 2 576 577
0 622 6 4 2 578 579
0 627 6 4 2 580 581
0 632 6 4 2 582 583
0 637 6 4 2 584 585
0 642 6 2 2 586 587
0 645 6 2 2 588 589
0 648 6 2 2 590 591
0 651 6 2 2 592 593
0 654 6 2 2 594 595
0 657 6 2 2 596 597
0 660 6 2 2 598 599
0 663 6 2 2 600 601
0 666 6 2 2 603 608
0 669 6 2 2 613 618
0 672 6 2 2 604 614
0 675 6 2 2 609 619
0 678 6 2 2 623 628
0 681 6 2 2 633 638
0 684 6 2 2 624 634
0 687 6 2 2 629 639
0 690 6 1 2 605 667
0 691 6 1 2 610 668
0 692 6 1 2 615 670
0 693 6 1 2 620 671
0 694 6 1 2 606 673
0 695 6 1 2 616 674
0 696 6 1 2 611 676
0 697 6 1 2 621 677
0 698 6 1 2 625 679
0 699 6 1 2 630 680
0 700 6 1 2 635 682
0 701 6 1 2 640 683
0 702 6 1 2 626 685
0 703 6 1 2 636 686
0 704 6 1 2 631 688
0 705 6 1 2 641 689
0 706 6 2 2 690 691
0 709 6 2 2 692 693
0 712 6 2 2 694 695
0 715 6 2 2 696 697
0 718 6 2 2 698 699
0 721 6 2 2 700 701
0 724 6 2 2 702 703
0 727 6 2 2 704 705
0 730 6 2 2 243 719
0 733 6 2 2 246 722
0 736 6 2 2 249 725
0 739 6 2 2 252 728
0 742 6 2 2 255 707
0 745 6 2 2 258 710
0 748 6 2 2 261 713
0 751 6 2 2 264 716
0 754 6 1 2 244 731
0 755 6 1 2 720 732
0 756 6 1 2 247 734
0 757 6 1 2 723 735
0 758 6 1 2 250 737
0 759 6 1 2 726 738
0 760 6 1 2 253 740
0 761 6 1 2 729 741
0 762 6 1 2 256 743
0 763 6 1 2 708 744
0 764 6 1 2 259 746
0 765 6 1 2 711 747
0 766 6 1 2 262 749
0 767 6 1 2 714 750
0 768 6 1 2 265 752
0 769 6 1 2 717 753
0 770 6 2 2 754 755
0 773 6 2 2 756 757
0 776 6 2 2 758 759
0 779 6 2 2 760 761
0 782 6 2 2 762 763
0 785 6 2 2 764 765
0 788 6 2 2 766 767
0 791 6 2 2 768 769
0 794 6 2 2 643 771
0 797 6 2 2 646 774
0 800 6 2 2 649 777
0 803 6 2 2 652 780
0 806 6 2 2 655 783
0 809 6 2 2 658 786
0 812 6 2 2 661 789
0 815 6 2 2 664 792
0 818 6 1 2 644 795
0 819 6 1 2 772 796
0 820 6 1 2 647 798
0 821 6 1 2 775 799
0 822 6 1 2 650 801
0 823 6 1 2 778 802
0 824 6 1 2 653 804
0 825 6 1 2 781 805
0 826 6 1 2 656 807
0 827 6 1 2 784 808
0 828 6 1 2 659 810
0 829 6 1 2 787 811
0 830 6 1 2 662 813
0 831 6 1 2 790 814
0 832 6 1 2 665 816
0 833 6 1 2 793 817
0 834 6 12 2 818 819
0 847 6 12 2 820 821
0 860 6 12 2 822 823
0 873 6 12 2 824 825
0 886 6 12 2 828 829
0 899 6 12 2 832 833
0 912 6 12 2 830 831
0 925 6 12 2 826 827
0 938 5 1 1 835
0 939 5 1 1 848
0 940 5 1 1 861
0 941 5 1 1 836
0 942 5 1 1 849
0 943 5 1 1 874
0 944 5 1 1 837
0 945 5 1 1 862
0 946 5 1 1 875
0 947 5 1 1 850
0 948 5 1 1 863
0 949 5 1 1 876
0 950 5 1 1 887
0 951 5 1 1 900
0 952 5 1 1 888
0 953 5 1 1 913
0 954 5 1 1 926
0 955 5 1 1 901
0 956 5 1 1 927
0 957 5 1 1 914
0 958 5 1 1 928
0 959 5 1 1 889
0 960 5 1 1 915
0 961 5 1 1 929
0 962 5 1 1 890
0 963 5 1 1 902
0 964 5 1 1 930
0 965 5 1 1 916
0 966 5 1 1 903
0 967 5 1 1 891
0 968 5 1 1 917
0 969 5 1 1 904
0 970 5 1 1 851
0 971 5 1 1 877
0 972 5 1 1 852
0 973 5 1 1 864
0 974 5 1 1 838
0 975 5 1 1 878
0 976 5 1 1 839
0 977 5 1 1 865
0 978 7 1 4 938 939 940 879
0 979 7 1 4 941 942 866 943
0 980 7 1 4 944 853 945 946
0 981 7 1 4 840 947 948 949
0 982 7 1 4 958 959 960 905
0 983 7 1 4 961 962 918 963
0 984 7 1 4 964 892 965 966
0 985 7 1 4 931 967 968 969
0 986 3 4 4 978 979 980 981
0 991 3 4 4 982 983 984 985
0 996 7 4 5 932 950 919 951 987
0 1001 7 4 5 933 952 953 906 988
0 1006 7 4 5 954 893 920 955 989
0 1011 7 4 5 956 894 957 907 990
0 1016 7 4 5 841 970 867 971 992
0 1021 7 4 5 842 972 973 880 993
0 1026 7 4 5 974 854 868 975 994
0 1031 7 4 5 976 855 977 881 995
0 1036 7 2 2 843 997
0 1039 7 2 2 856 998
0 1042 7 2 2 869 999
0 1045 7 2 2 882 1000
0 1048 7 2 2 844 1002
0 1051 7 2 2 857 1003
0 1054 7 2 2 870 1004
0 1057 7 2 2 883 1005
0 1060 7 2 2 845 1007
0 1063 7 2 2 858 1008
0 1066 7 2 2 871 1009
0 1069 7 2 2 884 1010
0 1072 7 2 2 846 1012
0 1075 7 2 2 859 1013
0 1078 7 2 2 872 1014
0 1081 7 2 2 885 1015
0 1084 7 2 2 934 1017
0 1087 7 2 2 895 1018
0 1090 7 2 2 921 1019
0 1093 7 2 2 908 1020
0 1096 7 2 2 935 1022
0 1099 7 2 2 896 1023
0 1102 7 2 2 922 1024
0 1105 7 2 2 909 1025
0 1108 7 2 2 936 1027
0 1111 7 2 2 897 1028
0 1114 7 2 2 923 1029
0 1117 7 2 2 910 1030
0 1120 7 2 2 937 1032
0 1123 7 2 2 898 1033
0 1126 7 2 2 924 1034
0 1129 7 2 2 911 1035
0 1132 6 2 2 6 1037
0 1135 6 2 2 13 1040
0 1138 6 2 2 20 1043
0 1141 6 2 2 27 1046
0 1144 6 2 2 34 1049
0 1147 6 2 2 41 1052
0 1150 6 2 2 48 1055
0 1153 6 2 2 55 1058
0 1156 6 2 2 62 1061
0 1159 6 2 2 69 1064
0 1162 6 2 2 76 1067
0 1165 6 2 2 83 1070
0 1168 6 2 2 90 1073
0 1171 6 2 2 97 1076
0 1174 6 2 2 104 1079
0 1177 6 2 2 111 1082
0 1180 6 2 2 118 1085
0 1183 6 2 2 125 1088
0 1186 6 2 2 132 1091
0 1189 6 2 2 139 1094
0 1192 6 2 2 146 1097
0 1195 6 2 2 153 1100
0 1198 6 2 2 160 1103
0 1201 6 2 2 167 1106
0 1204 6 2 2 174 1109
0 1207 6 2 2 181 1112
0 1210 6 2 2 188 1115
0 1213 6 2 2 195 1118
0 1216 6 2 2 202 1121
0 1219 6 2 2 209 1124
0 1222 6 2 2 216 1127
0 1225 6 2 2 223 1130
0 1228 6 1 2 7 1133
0 1229 6 1 2 1038 1134
0 1230 6 1 2 14 1136
0 1231 6 1 2 1041 1137
0 1232 6 1 2 21 1139
0 1233 6 1 2 1044 1140
0 1234 6 1 2 28 1142
0 1235 6 1 2 1047 1143
0 1236 6 1 2 35 1145
0 1237 6 1 2 1050 1146
0 1238 6 1 2 42 1148
0 1239 6 1 2 1053 1149
0 1240 6 1 2 49 1151
0 1241 6 1 2 1056 1152
0 1242 6 1 2 56 1154
0 1243 6 1 2 1059 1155
0 1244 6 1 2 63 1157
0 1245 6 1 2 1062 1158
0 1246 6 1 2 70 1160
0 1247 6 1 2 1065 1161
0 1248 6 1 2 77 1163
0 1249 6 1 2 1068 1164
0 1250 6 1 2 84 1166
0 1251 6 1 2 1071 1167
0 1252 6 1 2 91 1169
0 1253 6 1 2 1074 1170
0 1254 6 1 2 98 1172
0 1255 6 1 2 1077 1173
0 1256 6 1 2 105 1175
0 1257 6 1 2 1080 1176
0 1258 6 1 2 112 1178
0 1259 6 1 2 1083 1179
0 1260 6 1 2 119 1181
0 1261 6 1 2 1086 1182
0 1262 6 1 2 126 1184
0 1263 6 1 2 1089 1185
0 1264 6 1 2 133 1187
0 1265 6 1 2 1092 1188
0 1266 6 1 2 140 1190
0 1267 6 1 2 1095 1191
0 1268 6 1 2 147 1193
0 1269 6 1 2 1098 1194
0 1270 6 1 2 154 1196
0 1271 6 1 2 1101 1197
0 1272 6 1 2 161 1199
0 1273 6 1 2 1104 1200
0 1274 6 1 2 168 1202
0 1275 6 1 2 1107 1203
0 1276 6 1 2 175 1205
0 1277 6 1 2 1110 1206
0 1278 6 1 2 182 1208
0 1279 6 1 2 1113 1209
0 1280 6 1 2 189 1211
0 1281 6 1 2 1116 1212
0 1282 6 1 2 196 1214
0 1283 6 1 2 1119 1215
0 1284 6 1 2 203 1217
0 1285 6 1 2 1122 1218
0 1286 6 1 2 210 1220
0 1287 6 1 2 1125 1221
0 1288 6 1 2 217 1223
0 1289 6 1 2 1128 1224
0 1290 6 1 2 224 1226
0 1291 6 1 2 1131 1227
0 1292 6 1 2 1228 1229
0 1293 6 1 2 1230 1231
0 1294 6 1 2 1232 1233
0 1295 6 1 2 1234 1235
0 1296 6 1 2 1236 1237
0 1297 6 1 2 1238 1239
0 1298 6 1 2 1240 1241
0 1299 6 1 2 1242 1243
0 1300 6 1 2 1244 1245
0 1301 6 1 2 1246 1247
0 1302 6 1 2 1248 1249
0 1303 6 1 2 1250 1251
0 1304 6 1 2 1252 1253
0 1305 6 1 2 1254 1255
0 1306 6 1 2 1256 1257
0 1307 6 1 2 1258 1259
0 1308 6 1 2 1260 1261
0 1309 6 1 2 1262 1263
0 1310 6 1 2 1264 1265
0 1311 6 1 2 1266 1267
0 1312 6 1 2 1268 1269
0 1313 6 1 2 1270 1271
0 1314 6 1 2 1272 1273
0 1315 6 1 2 1274 1275
0 1316 6 1 2 1276 1277
0 1317 6 1 2 1278 1279
0 1318 6 1 2 1280 1281
0 1319 6 1 2 1282 1283
0 1320 6 1 2 1284 1285
0 1321 6 1 2 1286 1287
0 1322 6 1 2 1288 1289
0 1323 6 1 2 1290 1291
3 1324 9 0 1 1292
3 1325 9 0 1 1293
3 1326 9 0 1 1294
3 1327 9 0 1 1295
3 1328 9 0 1 1296
3 1329 9 0 1 1297
3 1330 9 0 1 1298
3 1331 9 0 1 1299
3 1332 9 0 1 1300
3 1333 9 0 1 1301
3 1334 9 0 1 1302
3 1335 9 0 1 1303
3 1336 9 0 1 1304
3 1337 9 0 1 1305
3 1338 9 0 1 1306
3 1339 9 0 1 1307
3 1340 9 0 1 1308
3 1341 9 0 1 1309
3 1342 9 0 1 1310
3 1343 9 0 1 1311
3 1344 9 0 1 1312
3 1345 9 0 1 1313
3 1346 9 0 1 1314
3 1347 9 0 1 1315
3 1348 9 0 1 1316
3 1349 9 0 1 1317
3 1350 9 0 1 1318
3 1351 9 0 1 1319
3 1352 9 0 1 1320
3 1353 9 0 1 1321
3 1354 9 0 1 1322
3 1355 9 0 1 1323
2 2 1 1
2 3 1 1
2 4 1 1
2 5 1 1
2 6 1 1
2 7 1 1
2 9 1 8
2 10 1 8
2 11 1 8
2 12 1 8
2 13 1 8
2 14 1 8
2 16 1 15
2 17 1 15
2 18 1 15
2 19 1 15
2 20 1 15
2 21 1 15
2 23 1 22
2 24 1 22
2 25 1 22
2 26 1 22
2 27 1 22
2 28 1 22
2 30 1 29
2 31 1 29
2 32 1 29
2 33 1 29
2 34 1 29
2 35 1 29
2 37 1 36
2 38 1 36
2 39 1 36
2 40 1 36
2 41 1 36
2 42 1 36
2 44 1 43
2 45 1 43
2 46 1 43
2 47 1 43
2 48 1 43
2 49 1 43
2 51 1 50
2 52 1 50
2 53 1 50
2 54 1 50
2 55 1 50
2 56 1 50
2 58 1 57
2 59 1 57
2 60 1 57
2 61 1 57
2 62 1 57
2 63 1 57
2 65 1 64
2 66 1 64
2 67 1 64
2 68 1 64
2 69 1 64
2 70 1 64
2 72 1 71
2 73 1 71
2 74 1 71
2 75 1 71
2 76 1 71
2 77 1 71
2 79 1 78
2 80 1 78
2 81 1 78
2 82 1 78
2 83 1 78
2 84 1 78
2 86 1 85
2 87 1 85
2 88 1 85
2 89 1 85
2 90 1 85
2 91 1 85
2 93 1 92
2 94 1 92
2 95 1 92
2 96 1 92
2 97 1 92
2 98 1 92
2 100 1 99
2 101 1 99
2 102 1 99
2 103 1 99
2 104 1 99
2 105 1 99
2 107 1 106
2 108 1 106
2 109 1 106
2 110 1 106
2 111 1 106
2 112 1 106
2 114 1 113
2 115 1 113
2 116 1 113
2 117 1 113
2 118 1 113
2 119 1 113
2 121 1 120
2 122 1 120
2 123 1 120
2 124 1 120
2 125 1 120
2 126 1 120
2 128 1 127
2 129 1 127
2 130 1 127
2 131 1 127
2 132 1 127
2 133 1 127
2 135 1 134
2 136 1 134
2 137 1 134
2 138 1 134
2 139 1 134
2 140 1 134
2 142 1 141
2 143 1 141
2 144 1 141
2 145 1 141
2 146 1 141
2 147 1 141
2 149 1 148
2 150 1 148
2 151 1 148
2 152 1 148
2 153 1 148
2 154 1 148
2 156 1 155
2 157 1 155
2 158 1 155
2 159 1 155
2 160 1 155
2 161 1 155
2 163 1 162
2 164 1 162
2 165 1 162
2 166 1 162
2 167 1 162
2 168 1 162
2 170 1 169
2 171 1 169
2 172 1 169
2 173 1 169
2 174 1 169
2 175 1 169
2 177 1 176
2 178 1 176
2 179 1 176
2 180 1 176
2 181 1 176
2 182 1 176
2 184 1 183
2 185 1 183
2 186 1 183
2 187 1 183
2 188 1 183
2 189 1 183
2 191 1 190
2 192 1 190
2 193 1 190
2 194 1 190
2 195 1 190
2 196 1 190
2 198 1 197
2 199 1 197
2 200 1 197
2 201 1 197
2 202 1 197
2 203 1 197
2 205 1 204
2 206 1 204
2 207 1 204
2 208 1 204
2 209 1 204
2 210 1 204
2 212 1 211
2 213 1 211
2 214 1 211
2 215 1 211
2 216 1 211
2 217 1 211
2 219 1 218
2 220 1 218
2 221 1 218
2 222 1 218
2 223 1 218
2 224 1 218
2 234 1 233
2 235 1 233
2 236 1 233
2 237 1 233
2 238 1 233
2 239 1 233
2 240 1 233
2 241 1 233
2 243 1 242
2 244 1 242
2 246 1 245
2 247 1 245
2 249 1 248
2 250 1 248
2 252 1 251
2 253 1 251
2 255 1 254
2 256 1 254
2 258 1 257
2 259 1 257
2 261 1 260
2 262 1 260
2 264 1 263
2 265 1 263
2 267 1 266
2 268 1 266
2 270 1 269
2 271 1 269
2 273 1 272
2 274 1 272
2 276 1 275
2 277 1 275
2 279 1 278
2 280 1 278
2 282 1 281
2 283 1 281
2 285 1 284
2 286 1 284
2 288 1 287
2 289 1 287
2 291 1 290
2 292 1 290
2 294 1 293
2 295 1 293
2 297 1 296
2 298 1 296
2 300 1 299
2 301 1 299
2 303 1 302
2 304 1 302
2 306 1 305
2 307 1 305
2 309 1 308
2 310 1 308
2 312 1 311
2 313 1 311
2 315 1 314
2 316 1 314
2 318 1 317
2 319 1 317
2 321 1 320
2 322 1 320
2 324 1 323
2 325 1 323
2 327 1 326
2 328 1 326
2 330 1 329
2 331 1 329
2 333 1 332
2 334 1 332
2 336 1 335
2 337 1 335
2 339 1 338
2 340 1 338
2 342 1 341
2 343 1 341
2 345 1 344
2 346 1 344
2 348 1 347
2 349 1 347
2 351 1 350
2 352 1 350
2 354 1 353
2 355 1 353
2 357 1 356
2 358 1 356
2 360 1 359
2 361 1 359
2 427 1 426
2 428 1 426
2 430 1 429
2 431 1 429
2 433 1 432
2 434 1 432
2 436 1 435
2 437 1 435
2 439 1 438
2 440 1 438
2 442 1 441
2 443 1 441
2 445 1 444
2 446 1 444
2 448 1 447
2 449 1 447
2 451 1 450
2 452 1 450
2 454 1 453
2 455 1 453
2 457 1 456
2 458 1 456
2 460 1 459
2 461 1 459
2 463 1 462
2 464 1 462
2 466 1 465
2 467 1 465
2 469 1 468
2 470 1 468
2 472 1 471
2 473 1 471
2 475 1 474
2 476 1 474
2 478 1 477
2 479 1 477
2 481 1 480
2 482 1 480
2 484 1 483
2 485 1 483
2 487 1 486
2 488 1 486
2 490 1 489
2 491 1 489
2 493 1 492
2 494 1 492
2 496 1 495
2 497 1 495
2 499 1 498
2 500 1 498
2 502 1 501
2 503 1 501
2 505 1 504
2 506 1 504
2 508 1 507
2 509 1 507
2 511 1 510
2 512 1 510
2 514 1 513
2 515 1 513
2 517 1 516
2 518 1 516
2 520 1 519
2 521 1 519
2 523 1 522
2 524 1 522
2 526 1 525
2 527 1 525
2 529 1 528
2 530 1 528
2 532 1 531
2 533 1 531
2 535 1 534
2 536 1 534
2 538 1 537
2 539 1 537
2 541 1 540
2 542 1 540
2 544 1 543
2 545 1 543
2 547 1 546
2 548 1 546
2 550 1 549
2 551 1 549
2 553 1 552
2 554 1 552
2 556 1 555
2 557 1 555
2 559 1 558
2 560 1 558
2 562 1 561
2 563 1 561
2 565 1 564
2 566 1 564
2 568 1 567
2 569 1 567
2 603 1 602
2 604 1 602
2 605 1 602
2 606 1 602
2 608 1 607
2 609 1 607
2 610 1 607
2 611 1 607
2 613 1 612
2 614 1 612
2 615 1 612
2 616 1 612
2 618 1 617
2 619 1 617
2 620 1 617
2 621 1 617
2 623 1 622
2 624 1 622
2 625 1 622
2 626 1 622
2 628 1 627
2 629 1 627
2 630 1 627
2 631 1 627
2 633 1 632
2 634 1 632
2 635 1 632
2 636 1 632
2 638 1 637
2 639 1 637
2 640 1 637
2 641 1 637
2 643 1 642
2 644 1 642
2 646 1 645
2 647 1 645
2 649 1 648
2 650 1 648
2 652 1 651
2 653 1 651
2 655 1 654
2 656 1 654
2 658 1 657
2 659 1 657
2 661 1 660
2 662 1 660
2 664 1 663
2 665 1 663
2 667 1 666
2 668 1 666
2 670 1 669
2 671 1 669
2 673 1 672
2 674 1 672
2 676 1 675
2 677 1 675
2 679 1 678
2 680 1 678
2 682 1 681
2 683 1 681
2 685 1 684
2 686 1 684
2 688 1 687
2 689 1 687
2 707 1 706
2 708 1 706
2 710 1 709
2 711 1 709
2 713 1 712
2 714 1 712
2 716 1 715
2 717 1 715
2 719 1 718
2 720 1 718
2 722 1 721
2 723 1 721
2 725 1 724
2 726 1 724
2 728 1 727
2 729 1 727
2 731 1 730
2 732 1 730
2 734 1 733
2 735 1 733
2 737 1 736
2 738 1 736
2 740 1 739
2 741 1 739
2 743 1 742
2 744 1 742
2 746 1 745
2 747 1 745
2 749 1 748
2 750 1 748
2 752 1 751
2 753 1 751
2 771 1 770
2 772 1 770
2 774 1 773
2 775 1 773
2 777 1 776
2 778 1 776
2 780 1 779
2 781 1 779
2 783 1 782
2 784 1 782
2 786 1 785
2 787 1 785
2 789 1 788
2 790 1 788
2 792 1 791
2 793 1 791
2 795 1 794
2 796 1 794
2 798 1 797
2 799 1 797
2 801 1 800
2 802 1 800
2 804 1 803
2 805 1 803
2 807 1 806
2 808 1 806
2 810 1 809
2 811 1 809
2 813 1 812
2 814 1 812
2 816 1 815
2 817 1 815
2 835 1 834
2 836 1 834
2 837 1 834
2 838 1 834
2 839 1 834
2 840 1 834
2 841 1 834
2 842 1 834
2 843 1 834
2 844 1 834
2 845 1 834
2 846 1 834
2 848 1 847
2 849 1 847
2 850 1 847
2 851 1 847
2 852 1 847
2 853 1 847
2 854 1 847
2 855 1 847
2 856 1 847
2 857 1 847
2 858 1 847
2 859 1 847
2 861 1 860
2 862 1 860
2 863 1 860
2 864 1 860
2 865 1 860
2 866 1 860
2 867 1 860
2 868 1 860
2 869 1 860
2 870 1 860
2 871 1 860
2 872 1 860
2 874 1 873
2 875 1 873
2 876 1 873
2 877 1 873
2 878 1 873
2 879 1 873
2 880 1 873
2 881 1 873
2 882 1 873
2 883 1 873
2 884 1 873
2 885 1 873
2 887 1 886
2 888 1 886
2 889 1 886
2 890 1 886
2 891 1 886
2 892 1 886
2 893 1 886
2 894 1 886
2 895 1 886
2 896 1 886
2 897 1 886
2 898 1 886
2 900 1 899
2 901 1 899
2 902 1 899
2 903 1 899
2 904 1 899
2 905 1 899
2 906 1 899
2 907 1 899
2 908 1 899
2 909 1 899
2 910 1 899
2 911 1 899
2 913 1 912
2 914 1 912
2 915 1 912
2 916 1 912
2 917 1 912
2 918 1 912
2 919 1 912
2 920 1 912
2 921 1 912
2 922 1 912
2 923 1 912
2 924 1 912
2 926 1 925
2 927 1 925
2 928 1 925
2 929 1 925
2 930 1 925
2 931 1 925
2 932 1 925
2 933 1 925
2 934 1 925
2 935 1 925
2 936 1 925
2 937 1 925
2 987 1 986
2 988 1 986
2 989 1 986
2 990 1 986
2 992 1 991
2 993 1 991
2 994 1 991
2 995 1 991
2 997 1 996
2 998 1 996
2 999 1 996
2 1000 1 996
2 1002 1 1001
2 1003 1 1001
2 1004 1 1001
2 1005 1 1001
2 1007 1 1006
2 1008 1 1006
2 1009 1 1006
2 1010 1 1006
2 1012 1 1011
2 1013 1 1011
2 1014 1 1011
2 1015 1 1011
2 1017 1 1016
2 1018 1 1016
2 1019 1 1016
2 1020 1 1016
2 1022 1 1021
2 1023 1 1021
2 1024 1 1021
2 1025 1 1021
2 1027 1 1026
2 1028 1 1026
2 1029 1 1026
2 1030 1 1026
2 1032 1 1031
2 1033 1 1031
2 1034 1 1031
2 1035 1 1031
2 1037 1 1036
2 1038 1 1036
2 1040 1 1039
2 1041 1 1039
2 1043 1 1042
2 1044 1 1042
2 1046 1 1045
2 1047 1 1045
2 1049 1 1048
2 1050 1 1048
2 1052 1 1051
2 1053 1 1051
2 1055 1 1054
2 1056 1 1054
2 1058 1 1057
2 1059 1 1057
2 1061 1 1060
2 1062 1 1060
2 1064 1 1063
2 1065 1 1063
2 1067 1 1066
2 1068 1 1066
2 1070 1 1069
2 1071 1 1069
2 1073 1 1072
2 1074 1 1072
2 1076 1 1075
2 1077 1 1075
2 1079 1 1078
2 1080 1 1078
2 1082 1 1081
2 1083 1 1081
2 1085 1 1084
2 1086 1 1084
2 1088 1 1087
2 1089 1 1087
2 1091 1 1090
2 1092 1 1090
2 1094 1 1093
2 1095 1 1093
2 1097 1 1096
2 1098 1 1096
2 1100 1 1099
2 1101 1 1099
2 1103 1 1102
2 1104 1 1102
2 1106 1 1105
2 1107 1 1105
2 1109 1 1108
2 1110 1 1108
2 1112 1 1111
2 1113 1 1111
2 1115 1 1114
2 1116 1 1114
2 1118 1 1117
2 1119 1 1117
2 1121 1 1120
2 1122 1 1120
2 1124 1 1123
2 1125 1 1123
2 1127 1 1126
2 1128 1 1126
2 1130 1 1129
2 1131 1 1129
2 1133 1 1132
2 1134 1 1132
2 1136 1 1135
2 1137 1 1135
2 1139 1 1138
2 1140 1 1138
2 1142 1 1141
2 1143 1 1141
2 1145 1 1144
2 1146 1 1144
2 1148 1 1147
2 1149 1 1147
2 1151 1 1150
2 1152 1 1150
2 1154 1 1153
2 1155 1 1153
2 1157 1 1156
2 1158 1 1156
2 1160 1 1159
2 1161 1 1159
2 1163 1 1162
2 1164 1 1162
2 1166 1 1165
2 1167 1 1165
2 1169 1 1168
2 1170 1 1168
2 1172 1 1171
2 1173 1 1171
2 1175 1 1174
2 1176 1 1174
2 1178 1 1177
2 1179 1 1177
2 1181 1 1180
2 1182 1 1180
2 1184 1 1183
2 1185 1 1183
2 1187 1 1186
2 1188 1 1186
2 1190 1 1189
2 1191 1 1189
2 1193 1 1192
2 1194 1 1192
2 1196 1 1195
2 1197 1 1195
2 1199 1 1198
2 1200 1 1198
2 1202 1 1201
2 1203 1 1201
2 1205 1 1204
2 1206 1 1204
2 1208 1 1207
2 1209 1 1207
2 1211 1 1210
2 1212 1 1210
2 1214 1 1213
2 1215 1 1213
2 1217 1 1216
2 1218 1 1216
2 1220 1 1219
2 1221 1 1219
2 1223 1 1222
2 1224 1 1222
2 1226 1 1225
2 1227 1 1225
