//# 8 inputs
//# 19 outputs
//# 6 D-type flipflops
//# 103 inverters
//# 550 gates (350 ANDs + 0 NANDs + 200 ORs + 0 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;

  wire NM,NCK;
  trireg NQ,M;

  nmos N7 (M,D,NCK);
  not P3 (NM,M);
  nmos N9 (NQ,NM,CK);
  not P5 (Q,NQ);
  not P1 (NCK,CK);

endmodule

module s1488(GND,VDD,CK,CLR,v0,v1,v13_D_10,v13_D_11,v13_D_12,v13_D_13,v13_D_14,
  v13_D_15,
  v13_D_16,v13_D_17,v13_D_18,v13_D_19,v13_D_20,v13_D_21,v13_D_22,v13_D_23,
  v13_D_24,v13_D_6,v13_D_7,v13_D_8,v13_D_9,v2,v3,v4,v5,v6);
input GND,VDD,CK,CLR,v6,v5,v4,v3,v2,v1,v0;
output v13_D_20,v13_D_21,v13_D_16,v13_D_22,v13_D_19,v13_D_18,v13_D_11,v13_D_23,
  v13_D_6,v13_D_15,v13_D_9,v13_D_10,v13_D_8,v13_D_24,v13_D_14,v13_D_7,v13_D_17,
  v13_D_12,v13_D_13;

  wire v12,v13_D_5C,v11,v13_D_4C,v10,v13_D_3C,v9,v13_D_2C,v8,v13_D_1C,v7,
    v13_D_0C,v0E,v1E,v2E,v3E,v4E,v5E,v6E,v7E,v8E,v9E,v10E,v11E,v12E,C208DE,
    C208D,II101,IIII518,C129DE,C129D,II114,C193D,C124DE,C124D,II143,IIII393,
    C108DE,C108D,C81DE,C81D,C83DE,C83D,II159,IIII344,C166DE,C166D,C104DE,C104D,
    C218DE,C218D,C131DE,C131D,C165DE,C165D,C220DE,C220D,C117DE,C117D,C194DE,
    C194D,C191DE,C191D,C141DE,C141D,C118DE,C118D,C70DE,C70D,C30DE,C30D,C144DE,
    C144D,C138DE,C138D,C157DE,C157D,C90DE,C90D,II246,C79D,C49DE,C49D,II294,
    IIII352,C150D,II373,IIII194,C97D,C180DE,C180D,II662,Av13_D_20B,II659,
    Av13_D_21B,C195DE,C195D,II674,Av13_D_16B,II656,Av13_D_22B,II665,Av13_D_19B,
    II668,Av13_D_18B,II689,Av13_D_11B,II653,Av13_D_23B,II704,Av13_D_6B,II677,
    Av13_D_15B,II695,Av13_D_9B,II692,Av13_D_10B,II698,Av13_D_8B,II650,
    Av13_D_24B,II680,Av13_D_14B,II722,Av13_D_0B,II701,Av13_D_7B,II713,
    Av13_D_3B,II719,Av13_D_1B,II707,Av13_D_5B,II710,Av13_D_4B,II671,Av13_D_17B,
    II716,Av13_D_2B,v13_D_0,v13_D_3,v13_D_1,II686,Av13_D_12B,v13_D_5,v13_D_4,
    v13_D_2,II683,Av13_D_13B,IIII533,IIII510,IIII389,IIII559,IIII546,IIII479,
    IIII380,IIII287,IIII516,IIII520,II329,IIII555,IIII537,IIII489,IIII461,
    IIII427,II254,IIII554,IIII528,IIII444,IIII442,II368,IIII534,IIII471,
    IIII464,IIII453,IIII430,IIII425,IIII167,IIII547,IIII524,II142,IIII508,
    IIII501,IIII492,IIII409,IIII357,IIII317,IIII170,IIII336,IIII560,IIII538,
    IIII506,IIII476,IIII466,IIII447,IIII417,IIII415,IIII412,IIII396,IIII372,
    IIII366,IIII333,IIII315,C155D,IIII251,IIII200,IIII189,IIII291,C142D,
    IIII392,IIII323,C127D,IIII381,IIII321,C33D,IIII378,IIII390,IIII350,IIII354,
    IIII399,IIII320,IIII349,IIII318,IIII486,IIII152,IIII329,IIII171,IIII175,
    IIII439,IIII403,IIII387,IIII369,IIII328,IIII310,IIII239,II642,IIII332,
    IIII306,IIII395,IIII347,IIII494,IIII299,IIII43,IIII365,C56D,IIII326,
    IIII500,IIII483,IIII478,IIII470,IIII468,IIII449,IIII296,IIII269,IIII259,
    IIII232,IIII513,C77D,IIII356,C50D,IIII335,IIII495,IIII420,IIII460,IIII435,
    IIII359,IIII338,IIII482,IIII452,IIII441,IIII498,IIII406,IIII191,IIII186,
    IIII134,C151D,IIII176,C145D,IIII497,IIII405,IIII463,IIII346,IIII485,
    IIII383,IIII219,IIII398,IIII341,IIII163,IIII109,C179D,IIII224,C163D,
    IIII503,IIII473,IIII456,IIII429,IIII419,IIII402,IIII386,IIII374,IIII205,
    IIII342,C159D,IIII438,IIII436,IIII433,IIII339,IIII272,IIII247,IIII243,
    IIII229,IIII226,IIII215,IIII202,IIII182,IIII179,IIII161,IIII148,IIII140,
    IIII136,C47D,IIII75,IIII111,C98D,IIII210,C120D,IIII375,C86D,IIII141,C170D,
    IIII79,IIII31,IIII514,IIII505,IIII491,IIII475,IIII450,IIII414,IIII384,
    IIII362,IIII293,IIII278,IIII256,IIII253,IIII250,IIII151,IIII363,C178D,
    IIII423,IIII302,IIII284,IIII131,IIII64,IIII360,C59D,IIII457,IIII446,
    IIII432,IIII377,IIII371,IIII368,IIII325,IIII314,IIII275,IIII157,C82D,
    IIII308,C111D,IIII208,C122D,IIII234,C167D,IIII35,IIII95,C76D,IIII282,C36D,
    IIII237,C221D,IIII177,C137D,IIII80,C192D,IIII305,IIII266,IIII212,IIII145,
    IIII203,C34D,IIII209,C119D,IIII199,C63D,IIII288,C203D,IIII206,IIII233,
    C168D,IIII128,C69D,IIII281,C29D,IIII285,C222D,IIII158,C84D,IIII227,C139D,
    IIII197,C158D,IIII248,C45D,IIII86,C54D,IIII91,C148D,IIII213,C57D,IIII276,
    C27D,IIII303,C172D,IIII263,C41D,IIII113,C93D,IIII114,IIII220,C51D,IIII240,
    C125D,IIII130,C60D,IIII267,C214D,C213D,IIII260,C78D,IIII222,C156D,IIII297,
    C209D,IIII101,C128D,IIII41,C96D,IIII34,C91D,IIII294,C211D,IIII174,C143D,
    IIII173,C146D,IIII273,C201D,IIII218,C44D,IIII192,IIII66,C100D,IIII82,C217D,
    IIII44,C106D,IIII104,C107D,IIII223,C160D,IIII257,C215D,IIII39,C103D,
    IIII230,C109D,IIII98,C87D,C200D,IIII40,C92D,IIII245,C185D,IIII65,IIII270,
    C55D,IIII300,C105D,IIII280,C26D,IIII311,C71D,IIII164,C133D,IIII156,C80D,
    IIII216,C189D,IIII254,C39D,IIII58,C75D,IIII106,C114D,IIII62,C95D,IIII262,
    C42D,IIII236,C219D,IIII242,C130D,IIII73,C31D,IIII188,C175D,IIII196,C161D,
    IIII149,C112D,IIII169,IIII183,C183D,IIII117,C35D,IIII120,C123D,IIII160,
    C65D,IIII166,C205D,IIII133,C152D,IIII142,C169D,IIII146,C223D,IIII92,C140D,
    IIII137,C46D,IIII126,C58D,IIII71,C28D,IIII180,C173D,IIII63,C99D,IIII119,
    C126D,IIII97,C88D,C210D,IIII185,IIII69,C202D,IIII153,C52D,II548,C199D,
    IIII124,C164D,C216D,IIII46,C110D,IIII54,C186D,IIII127,C73D,IIII103,C115D,
    IIII116,C37D,IIII129,C72D,IIII100,C134D,IIII96,C85D,IIII29,C190D,IIII154,
    C40D,IIII88,C43D,IIII83,C225D,IIII51,C132D,IIII49,C176D,IIII123,C162D,
    IIII105,C113D,IIII27,C184D,IIII93,C147D,IIII59,C67D,IIII68,C206D,C153D,
    IIII84,C224D,IIII89,C48D,IIII76,C174D,IIII108,C181D,IIII78,C196D,IIII72,
    C38D,IIII52,C135D,IIII36,C89D,IIII87,C53D,IIII45,C116D,IIII38,C102D,IIII32,
    C207D,IIII60,C74D,IIII48,C177D,IIII55,C187D,IIII28,C188D,II491,II497,II610,
    II542;

  dff DFF_0(CK,v12,v13_D_5C);
  dff DFF_1(CK,v11,v13_D_4C);
  dff DFF_2(CK,v10,v13_D_3C);
  dff DFF_3(CK,v9,v13_D_2C);
  dff DFF_4(CK,v8,v13_D_1C);
  dff DFF_5(CK,v7,v13_D_0C);
  not NOT_0(v0E,v0);
  not NOT_1(v1E,v1);
  not NOT_2(v2E,v2);
  not NOT_3(v3E,v3);
  not NOT_4(v4E,v4);
  not NOT_5(v5E,v5);
  not NOT_6(v6E,v6);
  not NOT_7(v7E,v7);
  not NOT_8(v8E,v8);
  not NOT_9(v9E,v9);
  not NOT_10(v10E,v10);
  not NOT_11(v11E,v11);
  not NOT_12(v12E,v12);
  not NOT_13(C208DE,C208D);
  not NOT_14(II101,v9);
  not NOT_15(IIII518,II101);
  not NOT_16(C129DE,C129D);
  not NOT_17(II114,v2);
  not NOT_18(C193D,II114);
  not NOT_19(C124DE,C124D);
  not NOT_20(II143,v10E);
  not NOT_21(IIII393,II143);
  not NOT_22(C108DE,C108D);
  not NOT_23(C81DE,C81D);
  not NOT_24(C83DE,C83D);
  not NOT_25(II159,C83D);
  not NOT_26(IIII344,II159);
  not NOT_27(C166DE,C166D);
  not NOT_28(C104DE,C104D);
  not NOT_29(C218DE,C218D);
  not NOT_30(C131DE,C131D);
  not NOT_31(C165DE,C165D);
  not NOT_32(C220DE,C220D);
  not NOT_33(C117DE,C117D);
  not NOT_34(C194DE,C194D);
  not NOT_35(C191DE,C191D);
  not NOT_36(C141DE,C141D);
  not NOT_37(C118DE,C118D);
  not NOT_38(C70DE,C70D);
  not NOT_39(C30DE,C30D);
  not NOT_40(C144DE,C144D);
  not NOT_41(C138DE,C138D);
  not NOT_42(C157DE,C157D);
  not NOT_43(C90DE,C90D);
  not NOT_44(II246,v11);
  not NOT_45(C79D,II246);
  not NOT_46(C49DE,C49D);
  not NOT_47(II294,IIII352);
  not NOT_48(C150D,II294);
  not NOT_49(II373,IIII194);
  not NOT_50(C97D,II373);
  not NOT_51(C180DE,C180D);
  not NOT_52(II662,Av13_D_20B);
  not NOT_53(v13_D_20,II662);
  not NOT_54(II659,Av13_D_21B);
  not NOT_55(C195DE,C195D);
  not NOT_56(II674,Av13_D_16B);
  not NOT_57(II656,Av13_D_22B);
  not NOT_58(v13_D_21,II659);
  not NOT_59(II665,Av13_D_19B);
  not NOT_60(v13_D_16,II674);
  not NOT_61(v13_D_22,II656);
  not NOT_62(II668,Av13_D_18B);
  not NOT_63(v13_D_19,II665);
  not NOT_64(II689,Av13_D_11B);
  not NOT_65(II653,Av13_D_23B);
  not NOT_66(II704,Av13_D_6B);
  not NOT_67(v13_D_18,II668);
  not NOT_68(II677,Av13_D_15B);
  not NOT_69(II695,Av13_D_9B);
  not NOT_70(v13_D_11,II689);
  not NOT_71(v13_D_23,II653);
  not NOT_72(II692,Av13_D_10B);
  not NOT_73(v13_D_6,II704);
  not NOT_74(II698,Av13_D_8B);
  not NOT_75(v13_D_15,II677);
  not NOT_76(v13_D_9,II695);
  not NOT_77(II650,Av13_D_24B);
  not NOT_78(v13_D_10,II692);
  not NOT_79(II680,Av13_D_14B);
  not NOT_80(v13_D_8,II698);
  not NOT_81(v13_D_24,II650);
  not NOT_82(II722,Av13_D_0B);
  not NOT_83(II701,Av13_D_7B);
  not NOT_84(II713,Av13_D_3B);
  not NOT_85(II719,Av13_D_1B);
  not NOT_86(II707,Av13_D_5B);
  not NOT_87(II710,Av13_D_4B);
  not NOT_88(v13_D_14,II680);
  not NOT_89(II671,Av13_D_17B);
  not NOT_90(II716,Av13_D_2B);
  not NOT_91(v13_D_0,II722);
  not NOT_92(v13_D_7,II701);
  not NOT_93(v13_D_3,II713);
  not NOT_94(v13_D_1,II719);
  not NOT_95(II686,Av13_D_12B);
  not NOT_96(v13_D_5,II707);
  not NOT_97(v13_D_4,II710);
  not NOT_98(v13_D_17,II671);
  not NOT_99(v13_D_2,II716);
  not NOT_100(v13_D_12,II686);
  not NOT_101(II683,Av13_D_13B);
  not NOT_102(v13_D_13,II683);
  and AND2_0(IIII533,v9,v10);
  and AND2_1(IIII510,v9,v10);
  and AND3_0(IIII389,v8,v9,v10);
  and AND2_2(IIII559,v8,v11);
  and AND2_3(IIII546,v0,v11);
  and AND2_4(IIII479,v0,v11);
  and AND2_5(IIII380,v2,v11);
  and AND2_6(IIII287,v9,v11);
  and AND2_7(IIII516,v1,v12);
  and AND2_8(IIII520,v3E,v6E);
  and AND3_1(II329,v3,v7E,v10);
  and AND3_2(IIII555,v0,v8E,v11);
  and AND4_0(IIII537,v6E,v7E,v8E,v12);
  and AND2_9(IIII489,v8E,v11);
  and AND3_3(IIII461,v8E,v9,v12);
  and AND3_4(IIII427,v8E,v9,v10);
  and AND4_1(II254,v1,v6,v7E,v8E);
  and AND3_5(IIII554,v2E,v8,v9E);
  and AND2_10(IIII528,v9E,v11);
  and AND2_11(IIII444,v3E,v9E);
  and AND3_6(IIII442,v7E,v8E,v9E);
  and AND3_7(II368,v7,v8,v9E);
  and AND2_12(IIII534,v8E,v10E);
  and AND3_8(IIII471,v1,v10E,v12);
  and AND3_9(IIII464,v8E,v10E,v11);
  and AND2_13(IIII453,v10E,v12);
  and AND3_10(IIII430,v1E,v9,v10E);
  and AND2_14(IIII425,v8E,v10E);
  and AND3_11(IIII167,v8,v11,C129D);
  and AND2_15(IIII547,v10,v11E);
  and AND2_16(IIII524,v6,v11E);
  and AND3_12(II142,v7E,v9,v11E);
  and AND2_17(IIII508,v9E,v11E);
  and AND2_18(IIII501,v8E,v11E);
  and AND2_19(IIII492,v10,v11E);
  and AND2_20(IIII409,v9,v11E);
  and AND2_21(IIII357,v10,v11E);
  and AND2_22(IIII317,v10,v11E);
  and AND2_23(IIII170,v10,v11E);
  and AND2_24(IIII352,v8,C124D);
  and AND2_25(IIII336,C124D,v12);
  and AND2_26(IIII560,v7E,v12E);
  and AND2_27(IIII538,v8,v12E);
  and AND4_2(IIII506,v7E,v9,v10E,v12E);
  and AND4_3(IIII476,v8E,v9,v11E,v12E);
  and AND3_13(IIII466,v8E,v11E,v12E);
  and AND4_4(IIII447,v8E,v9,v10E,v12E);
  and AND3_14(IIII417,v5E,v11E,v12E);
  and AND3_15(IIII415,v8E,v11E,v12E);
  and AND3_16(IIII412,v3,v10E,v12E);
  and AND2_28(IIII396,v10E,v12E);
  and AND2_29(IIII372,C129D,v12E);
  and AND4_5(IIII366,v8E,v9,v11E,v12E);
  and AND2_30(IIII333,v11E,v12E);
  and AND3_17(IIII315,C155D,v12E,C129D);
  and AND3_18(IIII251,v6E,v11E,v12E);
  and AND2_31(IIII200,v12E,C124D);
  and AND2_32(IIII189,v7,v12E);
  and AND2_33(IIII291,C142D,v11);
  and AND2_34(IIII392,C81D,v11E);
  and AND2_35(IIII323,v10E,C127D);
  and AND2_36(IIII381,C166D,v11E);
  and AND3_19(IIII321,C33D,v11E,v12E);
  and AND4_6(IIII378,C218D,v5E,v9,v12E);
  and AND2_37(IIII390,C220D,v10E);
  and AND2_38(IIII350,v11,C117D);
  and AND2_39(IIII354,C191D,v11);
  and AND2_40(IIII399,v8,C141D);
  and AND2_41(IIII320,v11,C141D);
  and AND2_42(IIII349,C118D,v11E);
  and AND2_43(IIII318,v11,C118D);
  and AND4_7(IIII486,v6E,v8E,v12,C129DE);
  and AND3_20(IIII152,v8,v12E,C129DE);
  and AND3_21(IIII329,v9,v12,C30D);
  and AND2_44(IIII171,v8,C193D);
  and AND2_45(IIII175,v9,C144D);
  and AND3_22(IIII439,v6,v12,C124DE);
  and AND4_8(IIII403,v9,v12E,C124DE,II254);
  and AND3_23(IIII387,v8E,v9E,C124DE);
  and AND2_46(IIII369,v9,C124DE);
  and AND3_24(IIII328,v3,v12E,C124DE);
  and AND4_9(IIII310,v6E,v9,v12E,C124DE);
  and AND3_25(IIII239,v9,v12,C124DE);
  and AND3_26(II642,v7E,v8E,C124DE);
  and AND2_47(IIII332,C138D,v9E);
  and AND2_48(IIII306,C129DE,C138D);
  and AND2_49(IIII395,C157D,v9E);
  and AND2_50(IIII347,C90D,v10E);
  and AND3_27(IIII494,v8E,v10,C108DE);
  and AND2_51(IIII299,v11E,C108DE);
  and AND3_28(IIII43,v8,v10,C108DE);
  and AND3_29(IIII365,C56D,v8,v11);
  and AND2_52(IIII326,C81DE,C129D);
  and AND3_30(IIII500,v8,v11,C83DE);
  and AND4_10(IIII483,v8E,v9E,v11E,C83DE);
  and AND2_53(IIII478,v10E,C83DE);
  and AND3_31(IIII470,v8,v12E,C83DE);
  and AND2_54(IIII468,v9,C83DE);
  and AND2_55(IIII449,C108DE,C83DE);
  and AND4_11(IIII296,v8E,v9E,C124DE,C83DE);
  and AND3_32(IIII269,v11E,C108DE,C83DE);
  and AND3_33(IIII259,v12E,C129DE,C83DE);
  and AND2_56(IIII232,C165D,C83DE);
  and AND3_34(IIII513,v12E,C166DE,II142);
  and AND3_35(IIII194,v3,v12,C77D);
  and AND2_57(IIII356,C50D,v10E);
  and AND2_58(IIII335,v12E,C218DE);
  and AND3_36(IIII495,v9,v11,C131DE);
  and AND3_37(IIII420,v2E,v7,C131DE);
  and AND3_38(IIII460,v2E,v12E,C165DE);
  and AND2_59(IIII435,v12,C165DE);
  and AND2_60(IIII359,v12E,C165DE);
  and AND2_61(IIII338,C108D,C165DE);
  and AND2_62(IIII482,v2,C220DE);
  and AND2_63(IIII452,v12E,C220DE);
  and AND2_64(IIII441,v11,C220DE);
  and AND2_65(IIII498,v8,C117DE);
  and AND3_39(IIII406,v8,v11,C117DE);
  and AND3_40(IIII191,v8,v11,C117DE);
  and AND3_41(IIII186,v8,v11,C117DE);
  and AND3_42(IIII134,v7E,v10,C151D);
  and AND2_66(IIII176,v10E,C145D);
  and AND3_43(IIII497,v8E,v9E,C194DE);
  and AND3_44(IIII405,v8E,v9E,C194DE);
  and AND2_67(IIII463,C165DE,C191DE);
  and AND2_68(IIII346,v12,C191DE);
  and AND3_45(IIII485,v6,C141DE,C220DE);
  and AND2_69(IIII383,C70D,C141DE);
  and AND2_70(IIII219,C49D,v9);
  and AND2_71(IIII398,v12E,C118DE);
  and AND2_72(IIII341,v11E,C118DE);
  and AND3_46(IIII163,v11E,v12E,C118DE);
  and AND4_12(IIII109,C179D,v2,v8,v11);
  and AND3_47(IIII224,C163D,v8E,v11);
  and AND2_73(IIII503,v9E,C30DE);
  and AND2_74(IIII473,v0E,C30DE);
  and AND2_75(IIII456,v9,C30DE);
  and AND2_76(IIII429,v9E,C30DE);
  and AND4_13(IIII419,v5E,v7E,v8E,C30DE);
  and AND3_48(IIII402,v8,v9E,C30DE);
  and AND4_14(IIII386,v0,C104D,v8,C30DE);
  and AND2_77(IIII374,v9E,C30DE);
  and AND2_78(IIII205,v8E,C30DE);
  and AND2_79(IIII342,C159D,v8E);
  and AND3_49(IIII438,v0,v10,C144DE);
  and AND3_50(IIII436,v8E,v9,C144DE);
  and AND2_80(IIII433,v10,C144DE);
  and AND2_81(IIII339,v8E,C144DE);
  and AND2_82(IIII272,v10E,C144DE);
  and AND2_83(IIII247,v10,C144DE);
  and AND3_51(IIII243,C131D,v9,C144DE);
  and AND3_52(IIII229,v9,v10,C144DE);
  and AND3_53(IIII226,v8E,v10E,C144DE);
  and AND3_54(IIII215,v1,v9,C144DE);
  and AND4_15(IIII202,v9E,C144DE,C83DE,C194DE);
  and AND3_55(IIII182,v8E,v10E,C144DE);
  and AND3_56(IIII179,v9,v10,C144DE);
  and AND2_84(IIII161,C144DE,C191D);
  and AND3_57(IIII148,v9,v10E,C144DE);
  and AND3_58(IIII140,v8E,v10E,C144DE);
  and AND2_85(IIII136,C47D,C144DE);
  and AND2_86(IIII75,C129DE,C144DE);
  and AND2_87(IIII111,C98D,v10E);
  and AND2_88(IIII210,v9,C120D);
  and AND2_89(IIII375,C86D,v10E);
  and AND2_90(IIII141,C170D,v8);
  and AND2_91(IIII79,v8,C170D);
  and AND3_59(IIII31,C108DE,C83DE,II642);
  and AND4_16(IIII514,v2,v7,v9E,C138DE);
  and AND4_17(IIII505,v7,v8,C138DE,C191DE);
  and AND2_92(IIII491,v10E,C138DE);
  and AND3_60(IIII475,v2E,v8,C138DE);
  and AND4_18(IIII450,v3,v8,C138DE,C104DE);
  and AND2_93(IIII414,v6,C138DE);
  and AND2_94(IIII384,v10E,C138DE);
  and AND2_95(IIII362,v8,C138DE);
  and AND4_19(Av13_D_20B,C138DE,C220DE,C104D,II329);
  and AND3_61(IIII293,C138DE,C118DE,II368);
  and AND2_96(IIII278,v10E,C138DE);
  and AND3_62(IIII256,v9,v10,C138DE);
  and AND3_63(IIII253,v1E,v10E,C138DE);
  and AND3_64(IIII250,C77D,v3,C138DE);
  and AND2_97(IIII151,v9,C138DE);
  and AND2_98(IIII363,v1E,C178D);
  and AND2_99(IIII423,v3E,C157DE);
  and AND2_100(IIII302,v11E,C157DE);
  and AND2_101(IIII284,v11E,C157DE);
  and AND3_65(IIII131,v9,v11E,C157DE);
  and AND2_102(IIII64,v11E,C157DE);
  and AND2_103(IIII360,v3E,C59D);
  and AND3_66(IIII457,v6,C124DE,C90DE);
  and AND2_104(IIII446,v11E,C90DE);
  and AND2_105(IIII432,v7,C90DE);
  and AND3_67(IIII377,v7,v10,C90DE);
  and AND2_106(IIII371,v10E,C90DE);
  and AND2_107(IIII368,C30D,C90DE);
  and AND2_108(IIII325,v10,C90DE);
  and AND2_109(IIII314,v10,C90DE);
  and AND3_68(IIII275,v7,v8,C90DE);
  and AND2_110(IIII157,C82D,v9E);
  and AND2_111(IIII308,C111D,C144DE);
  and AND2_112(IIII208,C122D,v11E);
  and AND2_113(IIII234,v8,C167D);
  and AND4_20(IIII35,C79D,v7,v9,v12E);
  and AND2_114(IIII95,C76D,C81DE);
  and AND2_115(IIII282,C36D,v12);
  and AND3_69(IIII237,v7,v12E,C221D);
  and AND2_116(IIII177,C137D,C127D);
  and AND3_70(IIII80,v7,v12E,C192D);
  and AND2_117(IIII305,v9,C49DE);
  and AND3_71(IIII266,v7,C49DE,C220DE);
  and AND2_118(IIII212,v9E,C49DE);
  and AND3_72(IIII145,C49DE,C166DE,C220DE);
  and AND2_119(IIII203,C34D,v9);
  and AND2_120(IIII209,v8,C119D);
  and AND2_121(IIII199,v9E,C63D);
  and AND2_122(IIII288,v7E,C203D);
  and AND2_123(IIII206,v7,C150D);
  and AND2_124(IIII233,C168D,v8E);
  and AND2_125(IIII128,v8,C69D);
  and AND2_126(IIII281,v3E,C29D);
  and AND2_127(IIII285,C222D,v10E);
  and AND2_128(IIII158,C84D,v10E);
  and AND3_73(IIII227,C139D,v8,v10);
  and AND3_74(IIII197,C158D,v7,v11E);
  and AND2_129(IIII248,C45D,v10E);
  and AND2_130(IIII86,C54D,C165DE);
  and AND2_131(IIII91,C148D,C131DE);
  and AND2_132(IIII213,C57D,v10E);
  and AND4_21(IIII276,C27D,v7E,v9,v12E);
  and AND2_133(IIII303,C172D,v12E);
  and AND3_75(IIII263,v7E,v11,C41D);
  and AND3_76(IIII113,v2E,v12E,C93D);
  and AND2_134(IIII114,v9,C97D);
  and AND2_135(IIII220,C51D,v12);
  and AND2_136(IIII240,C125D,v9E);
  and AND2_137(IIII130,C60D,C83D);
  and AND3_77(IIII267,C214D,v7E,v10E);
  and AND4_22(Av13_D_21B,C213D,v7E,v10E,v12E);
  and AND2_138(IIII260,v3E,C78D);
  and AND2_139(IIII222,C156D,C83DE);
  and AND3_78(IIII297,C209D,C208D,v11);
  and AND3_79(IIII101,C127D,C128D,v12E);
  and AND3_80(IIII41,v7,v12E,C96D);
  and AND2_140(IIII34,C91D,C165DE);
  and AND4_23(IIII294,C211D,v3,v7E,v11E);
  and AND2_141(IIII174,v8E,C143D);
  and AND2_142(IIII173,C146D,v11E);
  and AND2_143(IIII273,C201D,v8);
  and AND3_81(IIII218,v12E,C44D,C83DE);
  and AND3_82(IIII192,v8E,v9E,C44D);
  and AND3_83(IIII66,v8E,v12E,C100D);
  and AND3_84(IIII82,v0E,C217D,C108DE);
  and AND2_144(IIII44,v2E,C106D);
  and AND3_85(IIII104,v3,C107D,v12);
  and AND3_86(IIII223,v7E,C160D,v9E);
  and AND2_145(IIII257,C215D,v9E);
  and AND2_146(IIII39,C103D,v10E);
  and AND2_147(IIII230,C109D,v10E);
  and AND3_87(IIII98,v8E,v12,C87D);
  and AND3_88(Av13_D_16B,C200D,v8,v10);
  and AND2_148(IIII40,v2,C92D);
  and AND2_149(IIII245,C185D,v8E);
  and AND2_150(IIII65,v9,C185D);
  and AND2_151(IIII270,v1E,C55D);
  and AND2_152(IIII300,v0E,C105D);
  and AND2_153(IIII280,v1E,C26D);
  and AND2_154(IIII311,C71D,v9E);
  and AND2_155(IIII164,C133D,v8E);
  and AND2_156(IIII156,C80D,v9);
  and AND2_157(IIII216,C189D,v9E);
  and AND2_158(IIII254,C39D,v8E);
  and AND2_159(IIII58,C75D,C129DE);
  and AND2_160(IIII106,v8E,C114D);
  and AND2_161(IIII62,v6E,C95D);
  and AND2_162(IIII262,C42D,v8);
  and AND3_89(IIII236,v2E,v8,C219D);
  and AND2_163(IIII242,C130D,C165DE);
  and AND3_90(IIII73,v7,C31D,v8);
  and AND2_164(IIII188,C175D,v11);
  and AND2_165(IIII196,C161D,v11);
  and AND2_166(IIII149,C112D,v10);
  and AND2_167(IIII169,C195D,v8E);
  and AND2_168(IIII183,C183D,v8);
  and AND2_169(IIII117,v8E,C35D);
  and AND2_170(IIII120,v7E,C123D);
  and AND2_171(IIII160,v8,C65D);
  and AND2_172(IIII166,C205D,v10);
  and AND2_173(IIII133,C152D,v9);
  and AND2_174(IIII142,v7E,C169D);
  and AND3_91(IIII146,C223D,v8E,v9E);
  and AND2_175(IIII92,v7,C140D);
  and AND2_176(IIII137,v8,C46D);
  and AND2_177(IIII126,v2,C58D);
  and AND2_178(IIII71,v2E,C28D);
  and AND2_179(IIII180,C173D,v9E);
  and AND2_180(IIII63,v8,C99D);
  and AND2_181(IIII119,C126D,v8);
  and AND2_182(IIII97,C88D,v11E);
  and AND3_92(Av13_D_18B,C210D,v7E,v12E);
  and AND2_183(IIII185,v8E,C195DE);
  and AND2_184(IIII69,v7,C202D);
  and AND2_185(IIII153,C52D,v8E);
  and AND3_93(II548,C199D,v4,v5E);
  and AND2_186(IIII124,C164D,v12E);
  and AND3_94(Av13_D_23B,C216D,v7E,v8E);
  and AND2_187(IIII46,v7,C110D);
  and AND2_188(IIII54,C186D,v9E);
  and AND2_189(IIII127,C73D,v10E);
  and AND2_190(IIII103,C115D,v10);
  and AND2_191(IIII116,C37D,v9);
  and AND2_192(IIII129,v8E,C72D);
  and AND2_193(IIII100,C134D,v9E);
  and AND2_194(IIII96,v8,C85D);
  and AND2_195(IIII29,C190D,v10);
  and AND2_196(IIII154,v2,C40D);
  and AND2_197(IIII88,v2E,C43D);
  and AND2_198(IIII83,C225D,v11);
  and AND2_199(IIII51,C132D,v7);
  and AND2_200(IIII49,v8,C176D);
  and AND2_201(IIII123,v8,C162D);
  and AND2_202(IIII105,v8,C113D);
  and AND2_203(IIII27,C184D,v7);
  and AND2_204(IIII93,v7E,C147D);
  and AND2_205(IIII59,v7,C67D);
  and AND2_206(IIII68,C206D,v12E);
  and AND3_95(Av13_D_15B,v7E,v12E,II548);
  and AND2_207(Av13_D_9B,C153D,v12E);
  and AND2_208(IIII84,v7E,C224D);
  and AND2_209(IIII89,v7,C48D);
  and AND2_210(IIII76,v7E,C174D);
  and AND2_211(IIII108,C181D,C83DE);
  and AND2_212(IIII78,v7E,C196D);
  and AND2_213(IIII72,C38D,v7E);
  and AND2_214(IIII52,C135D,v7E);
  and AND2_215(IIII36,v7E,C89D);
  and AND2_216(IIII87,C53D,v7E);
  and AND2_217(IIII45,C116D,v7E);
  and AND2_218(IIII38,C102D,v7E);
  and AND2_219(IIII32,C207D,v2);
  and AND2_220(IIII60,v7E,C74D);
  and AND2_221(IIII48,C177D,v8E);
  and AND2_222(IIII55,C187D,v12E);
  and AND2_223(IIII28,v7E,C188D);
  and AND2_224(v13_D_0C,v13_D_0,CLR);
  and AND2_225(v13_D_3C,v13_D_3,CLR);
  and AND2_226(v13_D_1C,v13_D_1,CLR);
  and AND2_227(v13_D_5C,v13_D_5,CLR);
  and AND2_228(v13_D_4C,v13_D_4,CLR);
  and AND2_229(v13_D_2C,v13_D_2,CLR);
  or OR2_0(C208D,v5,v4);
  or OR2_1(C155D,v2,v7);
  or OR2_2(C129D,v9,v10);
  or OR2_3(C124D,v10,v11);
  or OR2_4(C142D,v0,v12);
  or OR2_5(C108D,v9,v12);
  or OR2_6(C81D,v2E,v12);
  or OR2_7(C83D,v4E,v5E);
  or OR2_8(C127D,v5E,v4);
  or OR2_9(C166D,v3E,v6E);
  or OR2_10(C33D,v6E,v10);
  or OR2_11(C104D,v1,v6E);
  or OR2_12(C218D,v7E,v10);
  or OR2_13(C131D,v8E,v10);
  or OR2_14(C165D,v8E,v11);
  or OR2_15(C220D,v8E,v9E);
  or OR2_16(C117D,v9E,v2);
  or OR2_17(C194D,v0,v10E);
  or OR2_18(C191D,v10E,v9);
  or OR2_19(C141D,v10E,v12);
  or OR2_20(C118D,v2E,v10E);
  or OR2_21(C70D,v0,v11E);
  or OR2_22(C30D,v10E,v11E);
  or OR2_23(C144D,v11E,v12);
  or OR2_24(C138D,v11E,v12E);
  or OR2_25(C157D,v10E,v12E);
  or OR2_26(C90D,v9,v12E);
  or OR2_27(C56D,v9,IIII516);
  or OR2_28(C77D,C104D,v0E);
  or OR2_29(C50D,IIII520,v11);
  or OR2_30(C151D,IIII554,IIII555);
  or OR2_31(C145D,IIII528,v12);
  or OR2_32(C47D,IIII533,IIII534);
  or OR2_33(C49D,C141D,v11);
  or OR2_34(C179D,v10,IIII518);
  or OR2_35(C163D,C129DE,IIII510);
  or OR2_36(C159D,IIII546,IIII547);
  or OR2_37(C98D,C144D,IIII444);
  or OR2_38(C120D,C144D,IIII425);
  or OR2_39(C86D,v9,IIII524);
  or OR2_40(C170D,C124DE,v9E);
  or OR2_41(C178D,IIII559,IIII560);
  or OR2_42(C59D,IIII537,IIII538);
  or OR2_43(C82D,IIII392,IIII393);
  or OR2_44(C111D,C83DE,v2);
  or OR2_45(C122D,v12,IIII323);
  or OR2_46(C167D,IIII380,IIII381);
  or OR2_47(C76D,C131DE,IIII427);
  or OR2_48(C36D,C165DE,v10E);
  or OR2_49(C221D,IIII389,IIII390);
  or OR2_50(C137D,C117DE,IIII489);
  or OR2_51(C180D,C194DE,v11E);
  or OR2_52(C192D,v8,IIII354);
  or OR2_53(C34D,IIII320,IIII321);
  or OR2_54(C119D,IIII349,IIII350);
  or OR2_55(C63D,IIII317,IIII318);
  or OR2_56(C203D,C70DE,IIII508);
  or OR2_57(C168D,C159D,v9);
  or OR2_58(C69D,IIII328,IIII329);
  or OR2_59(C29D,C138DE,IIII466);
  or OR2_60(C222D,C138DE,IIII417);
  or OR2_61(C84D,C138DE,IIII344);
  or OR2_62(C139D,IIII332,IIII333);
  or OR2_63(C158D,IIII395,IIII396);
  or OR2_64(C45D,C90DE,v11E);
  or OR2_65(C54D,C90DE,IIII412);
  or OR2_66(C148D,C90DE,IIII409);
  or OR2_67(C57D,IIII365,IIII366);
  or OR2_68(C27D,IIII500,IIII501);
  or OR2_69(C172D,IIII478,IIII479);
  or OR2_70(C41D,IIII470,IIII471);
  or OR2_71(C93D,C191DE,IIII468);
  or OR2_72(C51D,IIII356,IIII357);
  or OR2_73(C125D,IIII335,IIII336);
  or OR2_74(C60D,IIII494,IIII495);
  or OR2_75(C214D,IIII460,IIII461);
  or OR2_76(C213D,IIII482,IIII483);
  or OR2_77(C78D,IIII452,IIII453);
  or OR2_78(C156D,IIII441,IIII442);
  or OR2_79(C209D,IIII497,IIII498);
  or OR2_80(C128D,IIII405,IIII406);
  or OR2_81(C96D,IIII463,IIII464);
  or OR2_82(C91D,IIII346,IIII347);
  or OR2_83(C211D,IIII485,IIII486);
  or OR3_0(C143D,C49DE,v9,IIII291);
  or OR2_84(C146D,IIII398,IIII399);
  or OR2_85(C201D,IIII503,v12E);
  or OR2_86(C44D,IIII473,C124DE);
  or OR2_87(C100D,IIII429,IIII430);
  or OR2_88(C217D,IIII419,IIII420);
  or OR2_89(C106D,IIII402,IIII403);
  or OR2_90(C107D,IIII386,IIII387);
  or OR2_91(C160D,IIII341,IIII342);
  or OR2_92(C215D,IIII438,IIII439);
  or OR2_93(C103D,IIII435,IIII436);
  or OR2_94(C109D,IIII338,IIII339);
  or OR2_95(C87D,IIII374,IIII375);
  or OR2_96(C200D,IIII513,IIII514);
  or OR2_97(C92D,IIII505,IIII506);
  or OR2_98(C185D,IIII491,IIII492);
  or OR2_99(C55D,IIII475,IIII476);
  or OR2_100(C105D,IIII449,IIII450);
  or OR2_101(C26D,IIII414,IIII415);
  or OR2_102(C71D,IIII383,IIII384);
  or OR2_103(C133D,C49DE,IIII278);
  or OR2_104(C80D,IIII250,IIII251);
  or OR2_105(C189D,IIII362,IIII363);
  or OR2_106(C39D,IIII423,v9);
  or OR2_107(C75D,IIII359,IIII360);
  or OR2_108(C114D,IIII456,IIII457);
  or OR2_109(C95D,IIII446,IIII447);
  or OR2_110(C42D,IIII432,IIII433);
  or OR2_111(C219D,IIII377,IIII378);
  or OR2_112(C130D,IIII371,IIII372);
  or OR2_113(C31D,IIII368,IIII369);
  or OR2_114(C175D,IIII325,IIII326);
  or OR2_115(C161D,IIII314,IIII315);
  or OR2_116(C112D,IIII308,v9E);
  or OR2_117(C195D,C180DE,v9);
  or OR2_118(C183D,IIII305,IIII306);
  or OR2_119(C35D,IIII202,IIII203);
  or OR4_0(C123D,C157DE,IIII208,IIII209,IIII210);
  or OR2_120(C65D,IIII199,IIII200);
  or OR2_121(C205D,IIII287,IIII288);
  or OR2_122(C152D,IIII205,IIII206);
  or OR4_1(C169D,IIII232,IIII233,v12,IIII234);
  or OR2_123(C223D,IIII284,IIII285);
  or OR2_124(C140D,IIII226,IIII227);
  or OR2_125(C46D,IIII247,IIII248);
  or OR2_126(C58D,IIII212,IIII213);
  or OR2_127(C28D,IIII275,IIII276);
  or OR2_128(C173D,IIII302,IIII303);
  or OR3_1(C99D,IIII111,IIII113,IIII114);
  or OR2_129(C126D,IIII239,IIII240);
  or OR2_130(Av13_D_22B,IIII266,IIII267);
  or OR2_131(C88D,IIII259,IIII260);
  or OR2_132(C210D,IIII296,IIII297);
  or OR2_133(Av13_D_19B,IIII293,IIII294);
  or OR3_2(II491,IIII173,IIII174,IIII175);
  or OR2_134(C202D,IIII272,IIII273);
  or OR3_3(C52D,IIII218,IIII219,IIII220);
  or OR2_135(C199D,IIII191,IIII192);
  or OR3_4(C164D,IIII222,IIII223,IIII224);
  or OR2_136(C216D,IIII256,IIII257);
  or OR2_137(C110D,IIII229,IIII230);
  or OR2_138(C186D,C49DE,IIII245);
  or OR2_139(C73D,IIII269,IIII270);
  or OR2_140(C115D,IIII299,IIII300);
  or OR3_5(C37D,IIII280,IIII281,IIII282);
  or OR2_141(C72D,IIII310,IIII311);
  or OR2_142(C134D,IIII163,IIII164);
  or OR3_6(C85D,IIII156,IIII157,IIII158);
  or OR2_143(C190D,IIII215,IIII216);
  or OR2_144(C40D,IIII253,IIII254);
  or OR2_145(C43D,IIII262,IIII263);
  or OR2_146(C225D,IIII236,IIII237);
  or OR2_147(C132D,IIII242,IIII243);
  or OR2_148(C176D,IIII188,IIII189);
  or OR2_149(C162D,IIII196,IIII197);
  or OR2_150(C113D,IIII148,IIII149);
  or OR3_7(II497,C208DE,C83DE,IIII169);
  or OR2_151(C184D,IIII182,IIII183);
  or OR3_8(C147D,IIII176,IIII177,II491);
  or OR2_152(C67D,IIII160,IIII161);
  or OR2_153(C206D,IIII166,IIII167);
  or OR2_154(C153D,IIII133,IIII134);
  or OR3_9(Av13_D_11B,IIII140,IIII141,IIII142);
  or OR2_155(C224D,IIII145,IIII146);
  or OR2_156(C48D,IIII136,IIII137);
  or OR2_157(C174D,IIII179,IIII180);
  or OR3_10(II610,IIII62,IIII63,IIII64);
  or OR2_158(Av13_D_6B,IIII119,IIII120);
  or OR2_159(C181D,IIII185,IIII186);
  or OR4_2(C196D,IIII170,v12,IIII171,II497);
  or OR3_11(II542,IIII126,IIII127,IIII128);
  or OR2_160(C38D,IIII116,IIII117);
  or OR2_161(C135D,IIII100,IIII101);
  or OR4_3(C89D,IIII95,IIII96,IIII97,IIII98);
  or OR4_4(C53D,IIII151,IIII152,IIII153,IIII154);
  or OR2_162(Av13_D_10B,IIII123,IIII124);
  or OR4_5(C116D,IIII103,IIII104,IIII105,IIII106);
  or OR3_12(C102D,IIII65,IIII66,II610);
  or OR3_13(Av13_D_8B,IIII91,IIII92,IIII93);
  or OR2_163(C207D,IIII68,IIII69);
  or OR4_6(C74D,IIII129,IIII130,IIII131,II542);
  or OR3_14(Av13_D_24B,IIII82,IIII83,IIII84);
  or OR2_164(C177D,IIII75,IIII76);
  or OR2_165(C187D,IIII108,IIII109);
  or OR3_15(Av13_D_14B,IIII78,IIII79,IIII80);
  or OR3_16(Av13_D_0B,IIII71,IIII72,IIII73);
  or OR2_166(Av13_D_7B,IIII51,IIII52);
  or OR3_17(Av13_D_3B,IIII34,IIII35,IIII36);
  or OR4_7(Av13_D_1B,IIII86,IIII87,IIII88,IIII89);
  or OR4_8(Av13_D_5B,IIII43,IIII44,IIII45,IIII46);
  or OR4_9(Av13_D_4B,IIII38,IIII39,IIII40,IIII41);
  or OR2_167(Av13_D_17B,IIII31,IIII32);
  or OR3_18(Av13_D_2B,IIII58,IIII59,IIII60);
  or OR2_168(Av13_D_12B,IIII48,IIII49);
  or OR2_169(C188D,IIII54,IIII55);
  or OR3_19(Av13_D_13B,IIII27,IIII28,IIII29);

endmodule