1 0 0 5 0
1 1 0 5 0
1 2 0 6 0
1 3 0 6 0
1 4 0 6 0
1 5 0 6 0
1 6 0 6 0
1 7 0 4 0
1 8 0 6 0
1 9 0 6 0
1 10 0 5 0
1 11 0 4 0
1 12 0 6 0
1 13 0 5 0
1 14 0 6 0
1 15 0 6 0
1 16 0 5 0
1 17 0 6 0
1 18 0 6 0
1 19 0 5 0
1 20 0 6 0
1 21 0 6 0
1 22 0 5 0
1 23 0 5 0
1 24 0 6 0
1 25 0 5 0
1 26 0 6 0
1 27 0 5 0
1 28 0 6 0
1 29 0 5 0
1 30 0 6 0
1 31 0 5 0
1 32 0 1 0
1 33 0 1 0
1 34 0 1 0
1 35 0 1 0
1 36 0 1 0
1 37 0 1 0
1 38 0 1 0
1 39 0 1 0
1 40 0 8 0
2 41 1 0 
2 42 1 0 
2 43 1 0 
2 44 1 0 
2 45 1 0 
2 46 1 1 
2 47 1 1 
2 48 1 1 
2 49 1 1 
2 50 1 1 
2 51 1 2 
2 52 1 2 
2 53 1 2 
2 54 1 2 
2 55 1 2 
2 56 1 2 
2 57 1 3 
2 58 1 3 
2 59 1 3 
2 60 1 3 
2 61 1 3 
2 62 1 3 
2 63 1 4 
2 64 1 4 
2 65 1 4 
2 66 1 4 
2 67 1 4 
2 68 1 4 
2 69 1 5 
2 70 1 5 
2 71 1 5 
2 72 1 5 
2 73 1 5 
2 74 1 5 
2 75 1 6 
2 76 1 6 
2 77 1 6 
2 78 1 6 
2 79 1 6 
2 80 1 6 
2 81 1 7 
2 82 1 7 
2 83 1 7 
2 84 1 7 
2 85 1 8 
2 86 1 8 
2 87 1 8 
2 88 1 8 
2 89 1 8 
2 90 1 8 
2 91 1 9 
2 92 1 9 
2 93 1 9 
2 94 1 9 
2 95 1 9 
2 96 1 9 
2 97 1 10 
2 98 1 10 
2 99 1 10 
2 100 1 10 
2 101 1 10 
2 102 1 11 
2 103 1 11 
2 104 1 11 
2 105 1 11 
2 106 1 12 
2 107 1 12 
2 108 1 12 
2 109 1 12 
2 110 1 12 
2 111 1 12 
2 112 1 13 
2 113 1 13 
2 114 1 13 
2 115 1 13 
2 116 1 13 
2 117 1 14 
2 118 1 14 
2 119 1 14 
2 120 1 14 
2 121 1 14 
2 122 1 14 
2 123 1 15 
2 124 1 15 
2 125 1 15 
2 126 1 15 
2 127 1 15 
2 128 1 15 
2 129 1 16 
2 130 1 16 
2 131 1 16 
2 132 1 16 
2 133 1 16 
2 134 1 17 
2 135 1 17 
2 136 1 17 
2 137 1 17 
2 138 1 17 
2 139 1 17 
2 140 1 18 
2 141 1 18 
2 142 1 18 
2 143 1 18 
2 144 1 18 
2 145 1 18 
2 146 1 19 
2 147 1 19 
2 148 1 19 
2 149 1 19 
2 150 1 19 
2 151 1 20 
2 152 1 20 
2 153 1 20 
2 154 1 20 
2 155 1 20 
2 156 1 20 
2 157 1 21 
2 158 1 21 
2 159 1 21 
2 160 1 21 
2 161 1 21 
2 162 1 21 
2 163 1 22 
2 164 1 22 
2 165 1 22 
2 166 1 22 
2 167 1 22 
2 168 1 23 
2 169 1 23 
2 170 1 23 
2 171 1 23 
2 172 1 23 
2 173 1 24 
2 174 1 24 
2 175 1 24 
2 176 1 24 
2 177 1 24 
2 178 1 24 
2 179 1 25 
2 180 1 25 
2 181 1 25 
2 182 1 25 
2 183 1 25 
2 184 1 26 
2 185 1 26 
2 186 1 26 
2 187 1 26 
2 188 1 26 
2 189 1 26 
2 190 1 27 
2 191 1 27 
2 192 1 27 
2 193 1 27 
2 194 1 27 
2 195 1 28 
2 196 1 28 
2 197 1 28 
2 198 1 28 
2 199 1 28 
2 200 1 28 
2 201 1 29 
2 202 1 29 
2 203 1 29 
2 204 1 29 
2 205 1 29 
2 206 1 30 
2 207 1 30 
2 208 1 30 
2 209 1 30 
2 210 1 30 
2 211 1 30 
2 212 1 31 
2 213 1 31 
2 214 1 31 
2 215 1 31 
2 216 1 31 
2 217 1 40 
2 218 1 40 
2 219 1 40 
2 220 1 40 
2 221 1 40 
2 222 1 40 
2 223 1 40 
2 224 1 40 
0 225 6 2 2 32 217
0 226 6 3 2 34 218
0 227 6 3 2 35 219
0 228 6 3 2 33 220
0 229 6 2 2 38 221
0 230 5 3 1 210
0 231 5 2 1 167
0 232 5 3 1 188
0 233 5 3 1 145
0 234 5 2 1 49
0 235 5 2 1 133
0 236 5 3 1 199
0 237 5 3 1 178
0 238 5 4 1 45
0 239 5 3 1 156
0 240 5 3 1 61
0 241 5 3 1 56
0 242 6 2 2 36 222
0 243 5 3 1 105
0 244 5 3 1 162
0 245 6 2 2 37 223
0 246 5 3 1 89
0 247 5 4 1 183
0 248 5 2 1 100
0 249 5 3 1 139
0 250 5 4 1 205
0 251 5 4 1 216
0 252 5 3 1 83
0 253 5 2 1 172
0 254 5 3 1 73
0 255 5 3 1 80
0 256 6 3 2 39 224
0 257 5 4 1 194
0 258 5 4 1 150
0 259 5 3 1 67
0 260 5 3 1 111
0 261 5 4 1 115
0 262 5 3 1 128
2 263 1 225 
2 264 1 225 
2 265 1 226 
2 266 1 226 
2 267 1 226 
2 268 1 227 
2 269 1 227 
2 270 1 227 
2 271 1 228 
2 272 1 228 
2 273 1 228 
2 274 1 229 
2 275 1 229 
2 276 1 230 
2 277 1 230 
2 278 1 230 
2 279 1 231 
2 280 1 231 
2 281 1 232 
2 282 1 232 
2 283 1 232 
2 284 1 233 
2 285 1 233 
2 286 1 233 
2 287 1 234 
2 288 1 234 
2 289 1 235 
2 290 1 235 
2 291 1 236 
2 292 1 236 
2 293 1 236 
2 294 1 237 
2 295 1 237 
2 296 1 237 
2 297 1 238 
2 298 1 238 
2 299 1 238 
2 300 1 238 
2 301 1 239 
2 302 1 239 
2 303 1 239 
2 304 1 240 
2 305 1 240 
2 306 1 240 
2 307 1 241 
2 308 1 241 
2 309 1 241 
2 310 1 242 
2 311 1 242 
2 312 1 243 
2 313 1 243 
2 314 1 243 
2 315 1 244 
2 316 1 244 
2 317 1 244 
2 318 1 245 
2 319 1 245 
2 320 1 246 
2 321 1 246 
2 322 1 246 
2 323 1 247 
2 324 1 247 
2 325 1 247 
2 326 1 247 
2 327 1 248 
2 328 1 248 
2 329 1 249 
2 330 1 249 
2 331 1 249 
2 332 1 250 
2 333 1 250 
2 334 1 250 
2 335 1 250 
2 336 1 251 
2 337 1 251 
2 338 1 251 
2 339 1 251 
2 340 1 252 
2 341 1 252 
2 342 1 252 
2 343 1 253 
2 344 1 253 
2 345 1 254 
2 346 1 254 
2 347 1 254 
2 348 1 255 
2 349 1 255 
2 350 1 255 
2 351 1 256 
2 352 1 256 
2 353 1 256 
2 354 1 257 
2 355 1 257 
2 356 1 257 
2 357 1 257 
2 358 1 258 
2 359 1 258 
2 360 1 258 
2 361 1 258 
2 362 1 259 
2 363 1 259 
2 364 1 259 
2 365 1 260 
2 366 1 260 
2 367 1 260 
2 368 1 261 
2 369 1 261 
2 370 1 261 
2 371 1 261 
2 372 1 262 
2 373 1 262 
2 374 1 262 
0 375 6 1 2 159 358
0 376 6 1 2 148 315
0 377 6 1 2 170 279
0 378 6 1 2 165 343
0 379 4 1 2 160 359
0 380 4 1 2 149 316
0 381 6 1 2 142 289
0 382 6 1 2 131 284
0 383 5 2 1 266
0 384 6 1 2 175 307
0 385 6 1 2 53 294
0 386 4 1 2 77 281
0 387 4 1 2 186 348
0 388 6 1 2 78 282
0 389 6 1 2 187 349
0 390 4 1 2 176 308
0 391 4 1 2 54 295
0 392 5 2 1 269
0 393 6 1 2 153 304
0 394 6 1 2 59 301
0 395 4 1 2 203 291
0 396 4 1 2 197 332
0 397 6 1 2 204 292
0 398 6 1 2 198 333
0 399 4 1 2 154 305
0 400 4 1 2 60 302
0 401 6 1 2 181 271
0 402 4 1 2 182 272
0 403 5 2 1 273
0 404 6 1 2 71 336
0 405 6 1 2 214 345
0 406 4 1 2 208 354
0 407 4 1 2 192 276
0 408 6 1 2 209 355
0 409 6 1 2 193 277
0 410 4 1 2 72 337
0 411 4 1 2 215 346
0 412 6 1 2 143 320
0 413 6 1 2 87 285
0 414 6 1 2 104 327
0 415 6 1 2 99 312
0 416 6 1 2 93 274
0 417 3 1 2 94 275
0 418 6 1 2 166 278
0 419 6 1 2 211 280
0 420 6 1 2 48 283
0 421 6 1 2 189 287
0 422 4 1 2 144 321
0 423 4 1 2 88 286
0 424 6 1 2 132 288
0 425 6 1 2 50 290
0 426 6 1 2 177 293
0 427 6 1 2 200 296
0 428 6 1 2 155 362
0 429 6 1 2 65 303
0 430 6 1 2 55 306
0 431 6 1 2 62 309
0 432 6 1 2 161 372
0 433 6 1 2 125 317
0 434 6 1 2 119 318
0 435 3 1 2 120 319
0 436 6 1 2 108 322
0 437 6 1 2 90 365
0 438 6 1 2 138 328
0 439 6 1 2 101 331
0 440 3 1 2 95 368
0 441 6 1 2 96 369
0 442 6 1 2 171 342
0 443 6 1 2 84 344
0 444 6 1 2 79 347
0 445 6 1 2 74 350
0 446 5 2 1 352
0 447 3 1 2 121 360
0 448 6 1 2 122 361
0 449 6 1 2 126 370
0 450 6 1 2 114 373
0 451 4 1 2 109 363
0 452 4 1 2 66 366
0 453 6 1 2 110 364
0 454 6 1 2 68 367
0 455 4 1 2 127 371
0 456 4 1 2 116 374
0 457 6 1 2 376 375
0 458 6 2 2 378 377
0 459 4 1 2 380 379
0 460 6 4 2 382 381
0 461 6 1 2 385 384
0 462 4 1 2 387 386
0 463 6 1 2 389 388
0 464 4 1 2 391 390
0 465 6 1 2 394 393
0 466 4 1 2 396 395
0 467 6 1 2 398 397
0 468 4 1 2 400 399
0 469 6 1 2 405 404
0 470 4 1 2 407 406
0 471 6 1 2 409 408
0 472 4 1 2 411 410
0 473 6 1 2 413 412
0 474 6 2 2 415 414
0 475 7 2 2 417 416
0 476 6 4 2 419 418
0 477 6 4 2 421 420
0 478 4 1 2 423 422
0 479 6 2 2 425 424
0 480 6 5 2 427 426
0 481 6 2 2 429 428
0 482 6 3 2 431 430
0 483 6 2 2 433 432
0 484 6 2 2 435 434
0 485 6 2 2 437 436
0 486 6 2 2 439 438
0 487 6 2 2 441 440
0 488 6 2 2 443 442
0 489 6 5 2 445 444
0 490 6 2 2 448 447
0 491 6 1 2 450 449
0 492 4 1 2 452 451
0 493 6 1 2 454 453
0 494 4 1 2 456 455
2 495 1 383 
2 496 1 383 
2 497 1 392 
2 498 1 392 
2 499 1 403 
2 500 1 403 
2 501 1 446 
2 502 1 446 
0 503 6 1 2 462 461
0 504 6 1 2 464 463
0 505 6 1 2 466 465
0 506 6 1 2 468 467
0 507 6 1 2 499 323
0 508 4 1 2 500 324
0 509 6 1 2 470 469
0 510 6 1 2 472 471
0 511 6 1 2 492 491
0 512 6 1 2 494 493
2 513 1 458 
2 514 1 458 
2 515 1 460 
2 516 1 460 
2 517 1 460 
2 518 1 460 
2 519 1 474 
2 520 1 474 
2 521 1 475 
2 522 1 475 
2 523 1 476 
2 524 1 476 
2 525 1 476 
2 526 1 476 
2 527 1 477 
2 528 1 477 
2 529 1 477 
2 530 1 477 
2 531 1 479 
2 532 1 479 
2 533 1 480 
2 534 1 480 
2 535 1 480 
2 536 1 480 
2 537 1 480 
2 538 1 481 
2 539 1 481 
2 540 1 482 
2 541 1 482 
2 542 1 482 
2 543 1 483 
2 544 1 483 
2 545 1 484 
2 546 1 484 
2 547 1 485 
2 548 1 485 
2 549 1 486 
2 550 1 486 
2 551 1 487 
2 552 1 487 
2 553 1 488 
2 554 1 488 
2 555 1 489 
2 556 1 489 
2 557 1 489 
2 558 1 489 
2 559 1 489 
2 560 1 490 
2 561 1 490 
0 562 3 1 2 263 513
0 563 6 1 2 264 514
0 564 5 3 1 517
0 565 6 2 2 504 503
0 566 6 2 2 506 505
0 567 6 1 2 507 401
0 568 4 1 2 508 402
0 569 6 2 2 510 509
0 570 6 1 2 519 521
0 571 3 1 2 520 522
0 572 5 3 1 529
0 573 5 3 1 526
0 574 3 1 2 531 340
0 575 6 1 2 532 341
0 576 5 4 1 537
0 577 3 1 2 299 538
0 578 6 1 2 300 539
0 579 5 4 1 541
0 580 3 1 2 313 543
0 581 6 1 2 314 544
0 582 5 3 1 548
0 583 3 1 2 325 549
0 584 6 1 2 326 550
0 585 3 1 2 334 551
0 586 6 1 2 335 552
0 587 5 4 1 558
0 588 3 1 2 338 553
0 589 6 1 2 339 554
0 590 3 1 2 356 560
0 591 6 1 2 357 561
0 592 6 2 2 512 511
0 593 6 2 2 563 562
0 594 6 2 2 571 570
0 595 6 2 2 575 574
0 596 6 3 2 578 577
0 597 6 3 2 581 580
0 598 6 4 2 584 583
0 599 6 2 2 586 585
0 600 6 5 2 589 588
0 601 6 5 2 591 590
2 602 1 564 
2 603 1 564 
2 604 1 564 
2 605 1 565 
2 606 1 565 
2 607 1 566 
2 608 1 566 
2 609 1 569 
2 610 1 569 
2 611 1 572 
2 612 1 572 
2 613 1 572 
2 614 1 573 
2 615 1 573 
2 616 1 573 
2 617 1 576 
2 618 1 576 
2 619 1 576 
2 620 1 576 
2 621 1 579 
2 622 1 579 
2 623 1 579 
2 624 1 579 
2 625 1 582 
2 626 1 582 
2 627 1 582 
2 628 1 587 
2 629 1 587 
2 630 1 587 
2 631 1 587 
2 632 1 592 
2 633 1 592 
0 634 6 1 2 515 625
0 635 6 1 2 602 547
0 636 4 1 2 527 617
0 637 4 1 2 611 533
0 638 6 1 2 528 618
0 639 6 1 2 612 534
0 640 6 1 2 613 525
0 641 6 1 2 616 530
0 642 6 1 2 623 555
0 643 6 1 2 540 628
0 644 4 1 2 624 556
0 645 4 1 2 542 629
2 646 1 593 
2 647 1 593 
2 648 1 594 
2 649 1 594 
2 650 1 595 
2 651 1 595 
2 652 1 596 
2 653 1 596 
2 654 1 596 
2 655 1 597 
2 656 1 597 
2 657 1 597 
2 658 1 598 
2 659 1 598 
2 660 1 598 
2 661 1 598 
2 662 1 599 
2 663 1 599 
2 664 1 600 
2 665 1 600 
2 666 1 600 
2 667 1 600 
2 668 1 600 
2 669 1 601 
2 670 1 601 
2 671 1 601 
2 672 1 601 
2 673 1 601 
0 674 6 2 2 635 634
0 675 6 1 2 265 669
0 676 4 1 2 603 658
0 677 6 1 2 604 659
0 678 4 1 2 267 670
0 679 6 1 2 268 664
0 680 4 1 2 614 655
0 681 6 1 2 615 656
0 682 4 1 2 270 665
0 683 4 1 2 637 636
0 684 6 1 2 639 638
0 685 6 2 2 641 640
0 686 6 1 2 643 642
0 687 4 1 2 619 652
0 688 5 4 1 653
0 689 6 1 2 620 654
0 690 4 1 2 645 644
0 691 5 4 1 657
0 692 5 3 1 662
0 693 5 3 1 661
0 694 6 1 2 351 671
0 695 4 1 2 630 666
0 696 6 1 2 631 667
0 697 5 4 1 668
0 698 5 4 1 672
0 699 4 1 2 353 673
0 700 6 1 2 683 567
0 701 6 1 2 568 684
2 702 1 674 
2 703 1 674 
2 704 1 685 
2 705 1 685 
2 706 1 688 
2 707 1 688 
2 708 1 688 
2 709 1 688 
2 710 1 691 
2 711 1 691 
2 712 1 691 
2 713 1 691 
2 714 1 692 
2 715 1 692 
2 716 1 692 
2 717 1 693 
2 718 1 693 
2 719 1 693 
2 720 1 697 
2 721 1 697 
2 722 1 697 
2 723 1 697 
2 724 1 698 
2 725 1 698 
2 726 1 698 
2 727 1 698 
0 728 3 1 2 702 706
0 729 6 1 2 703 707
0 730 6 1 2 495 724
0 731 4 1 2 516 717
0 732 6 1 2 518 718
0 733 4 1 2 496 725
0 734 6 1 2 497 720
0 735 4 1 2 523 710
0 736 6 1 2 524 711
0 737 4 1 2 498 721
0 738 7 2 2 701 700
0 739 3 1 2 704 621
0 740 6 1 2 705 622
0 741 4 1 2 708 535
0 742 6 1 2 709 536
0 743 3 1 2 712 545
0 744 6 1 2 713 546
0 745 6 1 2 716 660
0 746 6 1 2 719 663
0 747 6 1 2 726 501
0 748 4 1 2 722 557
0 749 6 1 2 723 559
0 750 4 1 2 727 502
0 751 7 2 2 729 728
0 752 6 1 2 675 730
0 753 4 1 2 731 676
0 754 6 1 2 732 677
0 755 4 1 2 678 733
0 756 6 1 2 679 734
0 757 4 1 2 735 680
0 758 6 1 2 736 681
0 759 4 1 2 682 737
0 760 7 2 2 740 739
0 761 4 1 2 687 741
0 762 6 1 2 689 742
0 763 6 2 2 744 743
0 764 6 2 2 746 745
0 765 6 1 2 694 747
0 766 4 1 2 748 695
0 767 6 1 2 749 696
0 768 4 1 2 699 750
2 769 1 738 
2 770 1 738 
0 771 6 1 2 753 752
0 772 6 1 2 755 754
0 773 6 1 2 757 756
0 774 6 1 2 759 758
0 775 6 1 2 769 609
0 776 3 1 2 770 610
0 777 6 1 2 761 686
0 778 6 1 2 690 762
0 779 6 1 2 766 765
0 780 6 1 2 768 767
2 781 1 751 
2 782 1 751 
2 783 1 760 
2 784 1 760 
2 785 1 763 
2 786 1 763 
2 787 1 764 
2 788 1 764 
0 789 6 1 2 646 781
0 790 3 1 2 647 782
0 791 7 2 2 772 771
0 792 7 2 2 774 773
0 793 6 2 2 776 775
0 794 6 1 2 648 783
0 795 3 1 2 649 784
0 796 7 2 2 778 777
0 797 3 1 2 626 787
0 798 6 1 2 627 788
0 799 7 2 2 780 779
0 800 6 3 2 790 789
0 801 6 3 2 795 794
0 802 7 2 2 798 797
2 803 1 791 
2 804 1 791 
2 805 1 792 
2 806 1 792 
2 807 1 793 
2 808 1 793 
2 809 1 796 
2 810 1 796 
2 811 1 799 
2 812 1 799 
0 813 6 1 2 803 605
0 814 3 1 2 804 606
0 815 6 1 2 805 607
0 816 3 1 2 806 608
0 817 3 1 2 807 714
0 818 6 1 2 808 715
0 819 6 1 2 809 310
0 820 3 1 2 810 311
0 821 6 1 2 811 632
0 822 3 1 2 812 633
2 823 1 800 
2 824 1 800 
2 825 1 800 
2 826 1 801 
2 827 1 801 
2 828 1 801 
2 829 1 802 
2 830 1 802 
0 831 4 1 2 823 329
0 832 5 2 1 824
0 833 6 1 2 825 330
0 834 6 7 2 814 813
0 835 6 7 2 816 815
0 836 6 7 2 818 817
0 837 4 1 2 826 297
0 838 5 2 1 827
0 839 6 1 2 828 298
0 840 7 2 2 820 819
0 841 6 1 2 785 829
0 842 3 1 2 786 830
0 843 6 8 2 822 821
0 844 6 7 2 842 841
2 845 1 832 
2 846 1 832 
2 847 1 834 
2 848 1 834 
2 849 1 834 
2 850 1 834 
2 851 1 834 
2 852 1 834 
2 853 1 834 
2 854 1 835 
2 855 1 835 
2 856 1 835 
2 857 1 835 
2 858 1 835 
2 859 1 835 
2 860 1 835 
2 861 1 836 
2 862 1 836 
2 863 1 836 
2 864 1 836 
2 865 1 836 
2 866 1 836 
2 867 1 836 
2 868 1 838 
2 869 1 838 
2 870 1 840 
2 871 1 840 
2 872 1 843 
2 873 1 843 
2 874 1 843 
2 875 1 843 
2 876 1 843 
2 877 1 843 
2 878 1 843 
2 879 1 843 
0 880 4 1 2 847 861
0 881 5 2 1 876
0 882 4 1 2 136 845
0 883 6 1 2 137 846
0 884 5 3 1 859
0 885 5 2 1 866
0 886 5 4 1 853
0 887 4 3 2 860 867
0 888 4 1 2 43 868
0 889 6 1 2 44 869
0 890 6 1 2 650 870
0 891 3 1 2 651 871
2 892 1 844 
2 893 1 844 
2 894 1 844 
2 895 1 844 
2 896 1 844 
2 897 1 844 
2 898 1 844 
0 899 5 2 1 896
0 900 4 1 2 831 882
0 901 6 1 2 833 883
0 902 4 1 2 837 888
0 903 6 1 2 839 889
0 904 6 3 2 891 890
0 905 4 3 2 898 879
2 906 1 881 
2 907 1 881 
2 908 1 884 
2 909 1 884 
2 910 1 884 
2 911 1 885 
2 912 1 885 
2 913 1 886 
2 914 1 886 
2 915 1 886 
2 916 1 886 
2 917 1 887 
2 918 1 887 
2 919 1 887 
0 920 6 1 2 913 854
0 921 7 1 2 848 917
0 922 6 1 2 900 457
0 923 6 1 2 459 901
0 924 4 1 2 910 912
0 925 4 1 2 915 918
0 926 6 1 2 916 919
0 927 6 1 2 902 473
0 928 6 1 2 478 903
2 929 1 899 
2 930 1 899 
2 931 1 904 
2 932 1 904 
2 933 1 904 
2 934 1 905 
2 935 1 905 
2 936 1 905 
0 937 4 1 2 906 929
0 938 6 6 2 923 922
0 939 4 1 2 925 924
0 940 6 8 2 928 927
0 941 5 6 1 933
2 942 1 938 
2 943 1 938 
2 944 1 938 
2 945 1 938 
2 946 1 938 
2 947 1 938 
2 948 1 940 
2 949 1 940 
2 950 1 940 
2 951 1 940 
2 952 1 940 
2 953 1 940 
2 954 1 940 
2 955 1 940 
2 956 1 941 
2 957 1 941 
2 958 1 941 
2 959 1 941 
2 960 1 941 
2 961 1 941 
0 962 4 1 2 907 952
0 963 4 1 2 930 960
0 964 5 3 1 953
0 965 4 1 2 954 932
0 966 5 3 1 947
0 967 7 1 2 961 936
2 968 1 964 
2 969 1 964 
2 970 1 964 
2 971 1 966 
2 972 1 966 
2 973 1 966 
0 974 4 1 2 968 934
0 975 6 1 2 969 935
0 976 4 1 2 970 877
0 977 6 1 2 939 973
0 978 4 1 2 974 937
0 979 6 3 2 926 977
0 980 6 1 2 978 931
2 981 1 979 
2 982 1 979 
2 983 1 979 
0 984 6 2 2 975 980
0 985 7 2 2 963 981
0 986 6 1 2 982 878
0 987 7 1 2 983 955
0 988 4 1 2 986 897
0 989 7 4 2 967 987
2 990 1 984 
2 991 1 984 
2 992 1 985 
2 993 1 985 
0 994 6 1 2 990 942
0 995 5 2 1 991
0 996 7 4 2 962 992
0 997 7 4 2 976 993
0 998 7 4 2 965 988
2 999 1 989 
2 1000 1 989 
2 1001 1 989 
2 1002 1 989 
0 1003 4 1 2 994 909
0 1004 6 2 2 999 858
0 1005 6 2 2 1000 852
0 1006 6 2 2 1001 865
0 1007 6 2 2 1002 946
2 1008 1 995 
2 1009 1 995 
2 1010 1 996 
2 1011 1 996 
2 1012 1 996 
2 1013 1 996 
2 1014 1 997 
2 1015 1 997 
2 1016 1 997 
2 1017 1 997 
2 1018 1 998 
2 1019 1 998 
2 1020 1 998 
2 1021 1 998 
0 1022 4 1 2 1008 911
0 1023 7 4 2 880 1003
0 1024 4 1 2 1009 972
0 1025 6 2 2 1010 855
0 1026 6 2 2 1011 849
0 1027 6 2 2 1012 862
0 1028 6 2 2 1013 943
0 1029 6 2 2 1014 856
0 1030 6 2 2 1015 850
0 1031 6 2 2 1016 863
0 1032 6 2 2 1017 944
0 1033 6 2 2 1018 857
0 1034 6 2 2 1019 851
0 1035 6 2 2 1020 864
0 1036 6 2 2 1021 945
2 1037 1 1004 
2 1038 1 1004 
2 1039 1 1005 
2 1040 1 1005 
2 1041 1 1006 
2 1042 1 1006 
2 1043 1 1007 
2 1044 1 1007 
0 1045 6 2 2 1022 971
0 1046 7 4 2 921 1024
0 1047 6 1 2 57 1037
0 1048 3 1 2 58 1038
0 1049 6 1 2 51 1039
0 1050 3 1 2 52 1040
0 1051 6 1 2 46 1041
0 1052 3 1 2 47 1042
0 1053 6 1 2 41 1043
0 1054 3 1 2 42 1044
2 1055 1 1023 
2 1056 1 1023 
2 1057 1 1023 
2 1058 1 1023 
2 1059 1 1025 
2 1060 1 1025 
2 1061 1 1026 
2 1062 1 1026 
2 1063 1 1027 
2 1064 1 1027 
2 1065 1 1028 
2 1066 1 1028 
2 1067 1 1029 
2 1068 1 1029 
2 1069 1 1030 
2 1070 1 1030 
2 1071 1 1031 
2 1072 1 1031 
2 1073 1 1032 
2 1074 1 1032 
2 1075 1 1033 
2 1076 1 1033 
2 1077 1 1034 
2 1078 1 1034 
2 1079 1 1035 
2 1080 1 1035 
2 1081 1 1036 
2 1082 1 1036 
0 1083 6 2 2 1055 874
0 1084 6 2 2 1056 950
0 1085 6 2 2 1057 894
0 1086 6 2 2 1058 958
0 1087 6 1 2 123 1059
0 1088 3 1 2 124 1060
0 1089 6 1 2 117 1061
0 1090 3 1 2 118 1062
0 1091 6 1 2 112 1063
0 1092 3 1 2 113 1064
0 1093 6 1 2 106 1065
0 1094 3 1 2 107 1066
0 1095 6 1 2 102 1067
0 1096 3 1 2 103 1068
0 1097 6 1 2 97 1069
0 1098 3 1 2 98 1070
0 1099 6 1 2 91 1071
0 1100 3 1 2 92 1072
0 1101 6 1 2 85 1073
0 1102 3 1 2 86 1074
0 1103 6 1 2 81 1075
0 1104 3 1 2 82 1076
0 1105 6 1 2 75 1077
0 1106 3 1 2 76 1078
0 1107 6 1 2 69 1079
0 1108 3 1 2 70 1080
0 1109 6 1 2 63 1081
0 1110 3 1 2 64 1082
3 1111 6 0 2 1048 1047
3 1112 6 0 2 1050 1049
3 1113 6 0 2 1052 1051
3 1114 6 0 2 1054 1053
2 1115 1 1045 
2 1116 1 1045 
2 1117 1 1046 
2 1118 1 1046 
2 1119 1 1046 
2 1120 1 1046 
0 1121 4 4 2 920 1115
0 1122 4 1 2 1116 914
0 1123 6 2 2 1117 875
0 1124 6 2 2 1118 951
0 1125 6 2 2 1119 895
0 1126 6 2 2 1120 959
3 1127 6 0 2 1088 1087
3 1128 6 0 2 1090 1089
3 1129 6 0 2 1092 1091
3 1130 6 0 2 1094 1093
3 1131 6 0 2 1096 1095
3 1132 6 0 2 1098 1097
3 1133 6 0 2 1100 1099
3 1134 6 0 2 1102 1101
3 1135 6 0 2 1104 1103
3 1136 6 0 2 1106 1105
3 1137 6 0 2 1108 1107
3 1138 6 0 2 1110 1109
2 1139 1 1083 
2 1140 1 1083 
2 1141 1 1084 
2 1142 1 1084 
2 1143 1 1085 
2 1144 1 1085 
2 1145 1 1086 
2 1146 1 1086 
0 1147 7 4 2 1122 908
0 1148 6 1 2 168 1139
0 1149 3 1 2 169 1140
0 1150 6 1 2 163 1141
0 1151 3 1 2 164 1142
0 1152 6 1 2 157 1143
0 1153 3 1 2 158 1144
0 1154 6 1 2 151 1145
0 1155 3 1 2 152 1146
2 1156 1 1121 
2 1157 1 1121 
2 1158 1 1121 
2 1159 1 1121 
2 1160 1 1123 
2 1161 1 1123 
2 1162 1 1124 
2 1163 1 1124 
2 1164 1 1125 
2 1165 1 1125 
2 1166 1 1126 
2 1167 1 1126 
0 1168 6 2 2 1156 872
0 1169 6 2 2 1157 948
0 1170 6 2 2 1158 892
0 1171 6 2 2 1159 956
3 1172 6 0 2 1149 1148
3 1173 6 0 2 1151 1150
3 1174 6 0 2 1153 1152
3 1175 6 0 2 1155 1154
0 1176 6 1 2 146 1160
0 1177 3 1 2 147 1161
0 1178 6 1 2 140 1162
0 1179 3 1 2 141 1163
0 1180 6 1 2 134 1164
0 1181 3 1 2 135 1165
0 1182 6 1 2 129 1166
0 1183 3 1 2 130 1167
2 1184 1 1147 
2 1185 1 1147 
2 1186 1 1147 
2 1187 1 1147 
0 1188 6 2 2 1184 873
0 1189 6 2 2 1185 949
0 1190 6 2 2 1186 893
0 1191 6 2 2 1187 957
3 1192 6 0 2 1177 1176
3 1193 6 0 2 1179 1178
3 1194 6 0 2 1181 1180
3 1195 6 0 2 1183 1182
2 1196 1 1168 
2 1197 1 1168 
2 1198 1 1169 
2 1199 1 1169 
2 1200 1 1170 
2 1201 1 1170 
2 1202 1 1171 
2 1203 1 1171 
0 1204 6 1 2 212 1196
0 1205 3 1 2 213 1197
0 1206 6 1 2 206 1198
0 1207 3 1 2 207 1199
0 1208 6 1 2 201 1200
0 1209 3 1 2 202 1201
0 1210 6 1 2 195 1202
0 1211 3 1 2 196 1203
2 1212 1 1188 
2 1213 1 1188 
2 1214 1 1189 
2 1215 1 1189 
2 1216 1 1190 
2 1217 1 1190 
2 1218 1 1191 
2 1219 1 1191 
3 1220 6 0 2 1205 1204
3 1221 6 0 2 1207 1206
3 1222 6 0 2 1209 1208
3 1223 6 0 2 1211 1210
0 1224 6 1 2 190 1212
0 1225 3 1 2 191 1213
0 1226 6 1 2 184 1214
0 1227 3 1 2 185 1215
0 1228 6 1 2 179 1216
0 1229 3 1 2 180 1217
0 1230 6 1 2 173 1218
0 1231 3 1 2 174 1219
3 1232 6 0 2 1225 1224
3 1233 6 0 2 1227 1226
3 1234 6 0 2 1229 1228
3 1235 6 0 2 1231 1230
