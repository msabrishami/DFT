1    133    0    1    0
1    45    0    1    0
1    131    0    1    0
1    121    0    1    0
1    33    0    1    0
1    1    0    1    0
1    85    0    1    0
1    135    0    1    0
1    29    0    1    0
1    89    0    1    0
1    125    0    1    0
1    134    0    1    0
1    65    0    1    0
1    81    0    1    0
1    130    0    1    0
1    77    0    1    0
1    101    0    1    0
1    132    0    1    0
1    37    0    1    0
1    97    0    1    0
1    113    0    1    0
1    69    0    1    0
1    129    0    1    0
1    5    0    1    0
1    93    0    1    0
1    117    0    1    0
1    41    0    1    0
1    53    0    1    0
1    9    0    1    0
1    49    0    1    0
1    73    0    1    0
1    17    0    1    0
1    57    0    1    0
1    105    0    1    0
1    13    0    1    0
1    109    0    1    0
1    136    0    1    0
1    25    0    1    0
1    61    0    1    0
1    21    0    1    0
1    137    0    1    0
0    250    2    1    2    1    5
0    251    2    1    2    9    13
0    252    2    1    2    17    21
0    253    2    1    2    25    29
0    254    2    1    2    33    37
0    255    2    1    2    41    45
0    256    2    1    2    49    53
0    257    2    1    2    57    61
0    258    2    1    2    65    69
0    259    2    1    2    73    77
0    260    2    1    2    81    85
0    261    2    1    2    89    93
0    262    2    1    2    97    101
0    263    2    1    2    105    109
0    264    2    1    2    113    117
0    265    2    1    2    121    125
0    266    7    1    2    129    137
0    267    7    1    2    130    137
0    268    7    1    2    131    137
0    269    7    1    2    132    137
0    270    7    1    2    133    137
0    271    7    1    2    134    137
0    272    7    1    2    135    137
0    273    7    1    2    136    137
0    274    2    1    2    1    17
0    275    2    1    2    33    49
0    276    2    1    2    5    21
0    277    2    1    2    37    53
0    278    2    1    2    9    25
0    279    2    1    2    41    57
0    280    2    1    2    13    29
0    281    2    1    2    45    61
0    282    2    1    2    65    81
0    283    2    1    2    97    113
0    284    2    1    2    69    85
0    285    2    1    2    101    117
0    286    2    1    2    73    89
0    287    2    1    2    105    121
0    288    2    1    2    77    93
0    289    2    1    2    109    125
0    290    2    2    2    250    251
0    293    2    2    2    252    253
0    296    2    2    2    254    255
0    299    2    2    2    256    257
0    302    2    2    2    258    259
0    305    2    2    2    260    261
0    308    2    2    2    262    263
0    311    2    2    2    264    265
0    314    2    1    2    274    275
0    315    2    1    2    276    277
0    316    2    1    2    278    279
0    317    2    1    2    280    281
0    318    2    1    2    282    283
0    319    2    1    2    284    285
0    320    2    1    2    286    287
0    321    2    1    2    288    289
0    338    2    1    2    290    293
0    339    2    1    2    296    299
0    340    2    1    2    290    296
0    341    2    1    2    293    299
0    342    2    1    2    302    305
0    343    2    1    2    308    311
0    344    2    1    2    302    308
0    345    2    1    2    305    311
0    346    2    1    2    266    342
0    347    2    1    2    267    343
0    348    2    1    2    268    344
0    349    2    1    2    269    345
0    350    2    1    2    270    338
0    351    2    1    2    271    339
0    352    2    1    2    272    340
0    353    2    1    2    273    341
0    354    2    12    2    314    346
0    367    2    12    2    315    347
0    380    2    12    2    316    348
0    393    2    12    2    317    349
0    406    2    12    2    318    350
0    419    2    12    2    319    351
0    432    2    12    2    320    352
0    445    2    12    2    321    353
0    554    5    1    1    354
0    555    5    1    1    367
0    556    5    1    1    380
0    557    5    1    1    354
0    558    5    1    1    367
0    559    5    1    1    393
0    560    5    1    1    354
0    561    5    1    1    380
0    562    5    1    1    393
0    563    5    1    1    367
0    564    5    1    1    380
0    565    5    1    1    393
0    566    5    1    1    419
0    567    5    1    1    445
0    568    5    1    1    419
0    569    5    1    1    432
0    570    5    1    1    406
0    571    5    1    1    445
0    572    5    1    1    406
0    573    5    1    1    432
0    574    5    1    1    406
0    575    5    1    1    419
0    576    5    1    1    432
0    577    5    1    1    406
0    578    5    1    1    419
0    579    5    1    1    445
0    580    5    1    1    406
0    581    5    1    1    432
0    582    5    1    1    445
0    583    5    1    1    419
0    584    5    1    1    432
0    585    5    1    1    445
0    586    5    1    1    367
0    587    5    1    1    393
0    588    5    1    1    367
0    589    5    1    1    380
0    590    5    1    1    354
0    591    5    1    1    393
0    592    5    1    1    354
0    593    5    1    1    380
0    594    7    1    4    554    555    556    393
0    595    7    1    4    557    558    380    559
0    596    7    1    4    560    367    561    562
0    597    7    1    4    354    563    564    565
0    598    7    1    4    574    575    576    445
0    599    7    1    4    577    578    432    579
0    600    7    1    4    580    419    581    582
0    601    7    1    4    406    583    584    585
0    602    3    4    4    594    595    596    597
0    607    3    4    4    598    599    600    601
0    620    7    4    5    406    566    432    567    602
0    625    7    4    5    406    568    569    445    602
0    630    7    4    5    570    419    432    571    602
0    635    7    4    5    572    419    573    445    602
0    640    7    4    5    354    586    380    587    607
0    645    7    4    5    354    588    589    393    607
0    650    7    4    5    590    367    380    591    607
0    655    7    4    5    592    367    593    393    607
0    692    7    1    2    354    620
0    693    7    1    2    367    620
0    694    7    1    2    380    620
0    695    7    1    2    393    620
0    696    7    1    2    354    625
0    697    7    1    2    367    625
0    698    7    1    2    380    625
0    699    7    1    2    393    625
0    700    7    1    2    354    630
0    701    7    1    2    367    630
0    702    7    1    2    380    630
0    703    7    1    2    393    630
0    704    7    1    2    354    635
0    705    7    1    2    367    635
0    706    7    1    2    380    635
0    707    7    1    2    393    635
0    708    7    1    2    406    640
0    709    7    1    2    419    640
0    710    7    1    2    432    640
0    711    7    1    2    445    640
0    712    7    1    2    406    645
0    713    7    1    2    419    645
0    714    7    1    2    432    645
0    715    7    1    2    445    645
0    716    7    1    2    406    650
0    717    7    1    2    419    650
0    718    7    1    2    432    650
0    719    7    1    2    445    650
0    720    7    1    2    406    655
0    721    7    1    2    419    655
0    722    7    1    2    432    655
0    723    7    1    2    445    655
3    724    2    0    2    1    692
3    725    2    0    2    5    693
3    726    2    0    2    9    694
3    727    2    0    2    13    695
3    728    2    0    2    17    696
3    729    2    0    2    21    697
3    730    2    0    2    25    698
3    731    2    0    2    29    699
3    732    2    0    2    33    700
3    733    2    0    2    37    701
3    734    2    0    2    41    702
3    735    2    0    2    45    703
3    736    2    0    2    49    704
3    737    2    0    2    53    705
3    738    2    0    2    57    706
3    739    2    0    2    61    707
3    740    2    0    2    65    708
3    741    2    0    2    69    709
3    742    2    0    2    73    710
3    743    2    0    2    77    711
3    744    2    0    2    81    712
3    745    2    0    2    85    713
3    746    2    0    2    89    714
3    747    2    0    2    93    715
3    748    2    0    2    97    716
3    749    2    0    2    101    717
3    750    2    0    2    105    718
3    751    2    0    2    109    719
3    752    2    0    2    113    720
3    753    2    0    2    117    721
3    754    2    0    2    121    722
3    755    2    0    2    125    723
