1 1 0 2 0
1 4 0 6 0
1 11 0 2 0
1 14 0 2 0
1 17 0 2 0
1 20 0 2 0
1 23 0 1 0
1 24 0 1 0
1 25 0 1 0
1 26 0 1 0
1 27 0 3 0
1 31 0 2 0
1 34 0 2 0
1 37 0 2 0
1 40 0 2 0
1 43 0 2 0
1 46 0 2 0
1 49 0 2 0
1 52 0 1 0
1 53 0 1 0
1 54 0 6 0
1 61 0 2 0
1 64 0 2 0
1 67 0 2 0
1 70 0 2 0
1 73 0 2 0
1 76 0 2 0
1 79 0 1 0
1 80 0 1 0
1 81 0 1 0
1 82 0 1 0
1 83 0 2 0
1 86 0 1 0
1 87 0 1 0
1 88 0 2 0
1 91 0 2 0
1 94 0 2 0
1 97 0 2 0
1 100 0 2 0
1 103 0 2 0
1 106 0 2 0
1 109 0 2 0
1 112 0 1 0
1 113 0 1 0
1 114 0 1 0
1 115 0 1 0
1 116 0 1 0
1 117 0 1 0
1 118 0 1 0
1 119 0 1 0
1 120 0 1 0
1 121 0 1 0
1 122 0 1 0
1 123 0 2 0
1 126 0 1 0
1 127 0 1 0
1 128 0 1 0
1 129 0 1 0
1 130 0 1 0
1 131 0 1 0
1 132 0 2 0
1 135 0 1 0
1 136 0 1 0
1 137 0 2 0
1 140 0 1 0
1 141 0 3 0
1 145 0 1 0
1 146 0 2 0
1 149 0 2 0
1 152 0 2 0
1 155 0 2 0
1 158 0 2 0
1 161 0 2 0
1 164 0 2 0
1 167 0 2 0
1 170 0 2 0
1 173 0 2 0
1 176 0 2 0
1 179 0 2 0
1 182 0 2 0
1 185 0 2 0
1 188 0 2 0
1 191 0 2 0
1 194 0 2 0
1 197 0 2 0
1 200 0 2 0
1 203 0 2 0
1 206 0 2 0
1 209 0 1 0
1 210 0 6 0
1 217 0 1 0
1 218 0 6 0
1 225 0 1 0
1 226 0 6 0
1 233 0 1 0
1 234 0 6 0
1 241 0 1 0
1 242 0 2 0
1 245 0 2 0
1 248 0 2 0
1 251 0 2 0
1 254 0 2 0
1 257 0 6 0
1 264 0 1 0
1 265 0 6 0
1 272 0 1 0
1 273 0 6 0
1 280 0 1 0
1 281 0 6 0
1 288 0 1 0
1 289 0 2 0
1 292 0 1 0
1 293 0 5 0
1 299 0 2 0
1 302 0 4 0
1 307 0 1 0
1 308 0 6 0
1 315 0 1 0
1 316 0 6 0
1 323 0 1 0
1 324 0 6 0
1 331 0 1 0
1 332 0 2 0
1 335 0 2 0
1 338 0 2 0
1 341 0 6 0
1 348 0 2 0
1 351 0 6 0
1 358 0 2 0
1 361 0 4 0
1 366 0 2 0
1 369 0 2 0
1 372 0 1 0
1 373 0 1 0
1 374 0 11 0
1 386 0 2 0
1 389 0 10 0
1 400 0 10 0
1 411 0 10 0
1 422 0 12 0
1 435 0 10 0
1 446 0 10 0
1 457 0 10 0
1 468 0 10 0
1 479 0 10 0
1 490 0 12 0
1 503 0 10 0
1 514 0 8 0
1 523 0 10 0
1 534 0 10 0
1 545 0 3 0
1 549 0 2 0
1 552 0 3 0
1 556 0 2 0
1 559 0 2 0
1 562 0 3 0
1 566 0 4 0
1 571 0 2 0
1 574 0 2 0
1 577 0 2 0
1 580 0 2 0
1 583 0 4 0
1 588 0 2 0
1 591 0 1 0
1 592 0 2 0
1 595 0 1 0
1 596 0 1 0
1 597 0 1 0
1 598 0 1 0
1 599 0 3 0
1 603 0 3 0
1 607 0 2 0
1 610 0 2 0
1 613 0 2 0
1 616 0 2 0
1 619 0 5 0
1 625 0 5 0
1 631 0 1 0
3 709 9 0 1 142
3 816 9 0 1 294
0 1042 7 1 2 135 631
0 1043 5 1 1 591
3 1066 9 0 1 593
0 1067 5 12 1 595
0 1080 5 11 1 596
0 1092 5 11 1 597
0 1104 5 12 1 598
3 1137 5 0 1 546
3 1138 5 0 1 349
3 1139 5 0 1 367
3 1140 7 0 2 553 563
3 1141 5 0 1 550
3 1142 5 0 1 547
3 1143 5 0 1 548
3 1144 5 0 1 339
3 1145 5 0 1 359
0 1146 6 1 2 373 2
3 1147 7 0 2 143 145
0 1148 5 1 1 594
0 1149 5 1 1 1042
0 1150 7 1 2 1043 28
0 1151 7 1 2 387 557
3 1152 5 0 1 246
3 1153 5 0 1 554
3 1154 5 0 1 564
3 1155 5 0 1 560
0 1156 7 1 4 388 561 558 555
0 1157 5 3 1 567
0 1161 9 11 1 572
0 1173 9 11 1 575
0 1185 9 11 1 573
0 1197 9 11 1 576
0 1209 9 3 1 138
0 1213 9 2 1 139
0 1216 9 2 1 144
0 1219 5 3 1 584
0 1223 9 11 1 578
0 1235 9 11 1 581
0 1247 9 11 1 579
0 1259 9 11 1 582
0 1271 9 8 1 255
0 1280 9 11 1 252
0 1292 9 10 1 253
0 1303 9 11 1 249
0 1315 9 11 1 250
0 1327 9 11 1 611
0 1339 9 11 1 608
0 1351 9 11 1 614
0 1363 9 11 1 617
0 1375 9 2 1 211
0 1378 9 2 1 212
0 1381 9 2 1 219
0 1384 9 2 1 220
0 1387 9 2 1 227
0 1390 9 2 1 228
0 1393 9 2 1 235
0 1396 9 2 1 236
0 1415 9 2 1 258
0 1418 9 2 1 259
0 1421 9 2 1 266
0 1424 9 2 1 267
0 1427 9 2 1 274
0 1430 9 2 1 275
0 1433 9 2 1 282
0 1436 9 2 1 283
0 1455 9 6 1 336
0 1462 9 6 1 337
0 1469 9 5 1 207
0 1475 7 3 2 29 32
0 1479 9 2 1 3
0 1482 9 9 1 589
0 1492 9 2 1 295
0 1495 9 2 1 303
0 1498 9 2 1 309
0 1501 9 2 1 310
0 1504 9 2 1 317
0 1507 9 2 1 318
0 1510 9 2 1 325
0 1513 9 2 1 326
0 1516 9 2 1 342
0 1519 9 2 1 343
0 1522 9 2 1 352
0 1525 9 2 1 353
0 1542 9 2 1 260
0 1545 9 2 1 261
0 1548 9 2 1 268
0 1551 9 2 1 269
0 1554 9 2 1 276
0 1557 9 2 1 277
0 1560 9 2 1 284
0 1563 9 2 1 285
0 1566 9 6 1 333
0 1573 9 6 1 334
0 1580 9 2 1 551
0 1583 7 4 2 33 30
0 1588 5 5 1 590
0 1594 9 2 1 327
0 1597 9 2 1 328
0 1600 9 2 1 344
0 1603 9 2 1 345
0 1606 9 2 1 354
0 1609 9 2 1 355
0 1612 9 2 1 296
0 1615 9 2 1 304
0 1618 9 2 1 311
0 1621 9 2 1 312
0 1624 9 2 1 319
0 1627 9 2 1 320
0 1630 9 2 1 362
0 1633 9 2 1 363
0 1636 9 2 1 213
0 1639 9 2 1 214
0 1642 9 2 1 221
0 1645 9 2 1 222
0 1648 9 2 1 229
0 1651 9 2 1 230
0 1654 9 2 1 237
0 1657 9 2 1 238
0 1660 5 2 1 329
0 1663 9 11 1 243
0 1675 9 9 1 244
0 1685 9 11 1 256
0 1697 9 11 1 612
0 1709 9 11 1 609
0 1721 9 5 1 626
0 1727 9 3 1 620
0 1731 9 11 1 615
0 1743 9 11 1 618
0 1755 5 2 1 600
0 1758 5 2 1 604
0 1761 9 7 1 621
0 1769 9 7 1 627
0 1777 9 7 1 622
0 1785 9 7 1 628
0 1793 9 6 1 623
0 1800 9 6 1 629
0 1807 9 6 1 624
0 1814 9 6 1 630
0 1821 9 2 1 300
0 1824 9 2 1 447
0 1827 9 2 1 458
0 1830 9 2 1 469
0 1833 9 2 1 423
0 1836 9 2 1 436
0 1839 9 2 1 390
0 1842 9 2 1 401
0 1845 9 2 1 412
0 1848 9 2 1 375
0 1851 9 2 1 5
0 1854 9 2 1 448
0 1857 9 2 1 459
0 1860 9 2 1 470
0 1863 9 2 1 437
0 1866 9 2 1 391
0 1869 9 2 1 402
0 1872 9 2 1 413
0 1875 9 2 1 424
0 1878 9 2 1 376
0 1881 9 2 1 480
0 1884 9 2 1 491
0 1887 9 2 1 504
0 1890 9 2 1 515
0 1893 9 2 1 524
0 1896 9 2 1 535
0 1899 9 2 1 55
0 1902 9 2 1 481
0 1905 9 2 1 505
0 1908 9 2 1 516
0 1911 9 2 1 525
0 1914 9 2 1 536
0 1917 9 2 1 492
0 1920 9 2 1 364
0 1923 9 2 1 370
0 1926 9 2 1 346
0 1929 9 2 1 356
0 1932 9 2 1 313
0 1935 9 2 1 321
0 1938 9 2 1 297
0 1941 9 2 1 305
0 1944 9 2 1 286
0 1947 9 2 1 290
0 1950 9 2 1 270
0 1953 9 2 1 278
0 1956 9 2 1 239
0 1959 9 2 1 262
0 1962 9 2 1 223
0 1965 9 2 1 231
0 1968 9 2 1 215
3 1972 5 0 1 1146
3 2054 7 0 2 136 1148
3 2060 5 0 1 1150
3 2061 5 0 1 1151
3 2139 9 0 1 726
3 2142 9 0 1 731
3 2309 9 0 1 928
0 2349 7 1 2 666 517
0 2350 3 1 2 632 518
3 2387 9 0 1 991
3 2527 9 0 1 1224
3 2584 5 0 1 992
0 2585 7 1 3 171 681 692
0 2586 7 1 3 174 682 693
0 2587 7 1 3 168 683 694
0 2588 7 1 3 165 684 695
0 2589 7 1 3 162 685 696
3 2590 6 0 2 925 140
0 2591 7 1 3 186 703 715
0 2592 7 1 3 159 704 716
0 2593 7 1 3 153 705 717
0 2594 7 1 3 147 706 718
0 2595 7 1 3 172 736 747
0 2596 7 1 3 175 737 748
0 2597 7 1 3 169 738 749
0 2598 7 1 3 166 739 750
0 2599 7 1 3 163 740 751
0 2600 7 1 3 187 758 769
0 2601 7 1 3 160 759 770
0 2602 7 1 3 154 760 771
0 2603 7 1 3 148 761 772
0 2604 7 1 3 107 1116 1127
0 2605 7 1 3 62 832 843
0 2606 7 1 3 108 1084 1096
0 2607 7 1 3 50 1085 1097
0 2608 7 1 3 104 1086 1098
0 2609 7 1 3 41 1087 1099
0 2610 7 1 3 38 1088 1100
0 2611 7 1 3 21 833 844
0 2612 7 1 3 18 834 845
0 2613 7 1 3 71 835 846
0 2614 7 1 3 65 836 847
0 2615 7 1 3 51 1117 1128
0 2616 7 1 3 105 1118 1129
0 2617 7 1 3 42 1119 1130
0 2618 7 1 3 39 1120 1131
0 2619 7 1 3 22 854 865
0 2620 7 1 3 19 855 866
0 2621 7 1 3 72 856 867
0 2622 7 1 3 66 857 868
3 2623 5 0 1 926
0 2624 7 1 3 124 1162 601
0 2625 7 1 2 1179 1187
0 2626 7 1 3 63 858 869
0 2627 7 1 2 1164 1171
0 2628 5 1 1 1226
0 2629 5 1 1 1228
0 2630 5 1 1 1230
0 2631 5 1 1 1232
0 2632 5 1 1 1234
0 2633 5 1 1 1237
0 2634 5 1 1 1239
0 2635 5 1 1 1241
0 2636 5 1 1 1243
0 2637 5 1 1 1245
0 2638 5 1 1 1248
0 2639 5 1 1 1250
0 2640 5 1 1 1252
0 2641 5 1 1 1254
0 2642 5 1 1 1256
0 2643 5 1 1 1258
0 2644 5 1 1 1261
0 2645 5 1 1 1263
0 2646 5 1 1 1265
0 2647 9 5 1 727
0 2653 5 10 1 686
0 2664 5 10 1 697
0 2675 9 5 1 728
0 2681 5 10 1 707
0 2692 5 10 1 719
0 2703 7 1 3 180 708 720
0 2704 9 4 1 929
0 2709 5 1 1 1267
0 2710 5 1 1 1269
0 2711 5 1 1 1272
0 2712 5 1 1 1274
0 2713 5 1 1 1276
0 2714 5 1 1 1278
0 2715 5 1 1 1281
0 2716 5 1 1 1283
0 2717 5 1 1 1285
0 2718 5 1 1 1287
0 2719 5 1 1 1289
0 2720 5 1 1 1291
0 2721 5 1 1 1294
0 2722 9 5 1 729
0 2728 5 10 1 741
0 2739 5 10 1 752
0 2750 9 5 1 730
0 2756 5 10 1 762
0 2767 5 10 1 773
0 2778 7 1 3 181 763 774
0 2779 5 10 1 837
0 2790 5 10 1 848
0 2801 5 10 1 859
0 2812 5 10 1 870
0 2823 5 1 1 876
0 2824 5 1 1 878
0 2825 5 1 1 880
0 2826 5 1 1 882
0 2827 5 1 1 884
0 2828 5 1 1 886
0 2829 5 1 1 888
0 2830 5 1 1 890
0 2831 7 1 3 667 460 879
0 2832 7 1 3 668 471 883
0 2833 7 1 3 669 425 887
0 2834 7 1 3 670 438 891
0 2835 7 1 2 633 877
0 2836 7 1 2 634 881
0 2837 7 1 2 635 885
0 2838 7 1 2 636 889
0 2839 5 1 1 892
0 2840 5 1 1 894
0 2841 5 1 1 896
0 2842 5 1 1 898
0 2843 5 1 1 900
0 2844 5 1 1 902
0 2845 5 1 1 904
0 2846 5 1 1 906
0 2847 7 1 3 671 392 895
0 2848 7 1 3 672 403 899
0 2849 7 1 3 673 414 903
0 2850 7 1 3 674 377 907
0 2851 7 1 2 637 893
0 2852 7 1 2 638 897
0 2853 7 1 2 639 901
0 2854 7 1 2 640 905
0 2855 5 5 1 908
0 2861 5 5 1 914
0 2867 7 1 2 292 909
0 2868 7 1 2 288 910
0 2869 7 1 2 280 911
0 2870 7 1 2 272 912
0 2871 7 1 2 264 913
0 2872 7 1 2 241 915
0 2873 7 1 2 233 916
0 2874 7 1 2 225 917
0 2875 7 1 2 217 918
0 2876 7 1 2 209 919
0 2877 9 4 1 732
0 2882 5 8 1 930
0 2891 5 9 1 927
0 2901 5 1 1 939
0 2902 5 1 1 941
0 2903 5 1 1 943
0 2904 5 1 1 945
0 2905 5 1 1 947
0 2906 5 1 1 949
0 2907 7 1 2 809 942
0 2908 7 1 3 810 482 946
0 2909 7 1 3 811 493 950
0 2910 7 1 2 1050 940
0 2911 7 1 2 1051 944
0 2912 7 1 2 1052 948
0 2913 5 1 1 951
0 2914 5 1 1 953
0 2915 5 1 1 955
0 2916 5 1 1 957
0 2917 5 1 1 959
0 2918 5 1 1 961
0 2919 7 1 3 675 506 954
0 2920 5 1 1 2349
0 2921 7 1 3 676 526 958
0 2922 7 1 3 677 537 962
0 2923 7 1 2 641 952
0 2924 7 1 2 642 956
0 2925 7 1 2 643 960
0 2926 5 1 1 963
0 2927 5 1 1 965
0 2928 5 1 1 967
0 2929 5 1 1 969
0 2930 5 1 1 971
0 2931 5 1 1 973
0 2932 5 1 1 975
0 2933 5 1 1 977
0 2934 7 1 3 812 393 966
0 2935 7 1 3 813 404 970
0 2936 7 1 3 814 415 974
0 2937 7 1 3 815 378 978
0 2938 7 1 2 1053 964
0 2939 7 1 2 1054 968
0 2940 7 1 2 1055 972
0 2941 7 1 2 1056 976
0 2942 5 5 1 979
0 2948 5 5 1 985
0 2954 7 1 2 372 980
0 2955 7 1 2 368 981
0 2956 7 1 2 360 982
0 2957 7 1 2 350 983
0 2958 7 1 2 340 984
0 2959 7 1 2 331 986
0 2960 7 1 2 323 987
0 2961 7 1 2 315 988
0 2962 7 1 2 307 989
0 2963 7 1 2 301 990
0 2964 5 4 1 997
0 2969 7 1 2 84 998
0 2970 7 1 2 86 999
0 2971 7 1 2 89 1000
0 2972 7 1 2 90 1001
0 2973 5 1 1 1002
0 2974 5 1 1 1004
0 2975 5 1 1 1006
0 2976 5 1 1 1008
0 2977 5 1 1 1010
0 2978 5 1 1 1012
0 2979 7 1 3 821 507 1005
0 2980 7 1 2 822 519
0 2981 7 1 3 823 527 1009
0 2982 7 1 3 824 538 1013
0 2983 7 1 2 1061 1003
0 2984 3 1 2 1062 520
0 2985 7 1 2 1063 1007
0 2986 7 1 2 1064 1011
0 2987 5 1 1 1014
0 2988 5 1 1 1016
0 2989 5 1 1 1018
0 2990 5 1 1 1020
0 2991 5 1 1 1022
0 2992 5 1 1 1024
0 2993 7 1 2 825 1017
0 2994 7 1 3 826 483 1021
0 2995 7 1 3 827 494 1025
0 2996 7 1 2 1065 1015
0 2997 7 1 2 1068 1019
0 2998 7 1 2 1069 1023
0 2999 5 1 1 1026
0 3000 9 2 1 920
0 3003 9 2 1 921
0 3006 5 1 1 1028
0 3007 9 2 1 922
0 3010 9 2 1 923
0 3013 7 1 2 828 1027
0 3014 7 1 2 829 1029
0 3015 5 1 1 1030
0 3016 5 1 1 1032
0 3017 5 1 1 1034
0 3018 5 1 1 1036
0 3019 5 1 1 1038
0 3020 5 1 1 1040
0 3021 5 1 1 1044
0 3022 5 1 1 1046
0 3023 7 1 3 817 461 1033
0 3024 7 1 3 818 472 1037
0 3025 7 1 3 819 426 1041
0 3026 7 1 3 820 439 1047
0 3027 7 1 2 1057 1031
0 3028 7 1 2 1058 1035
0 3029 7 1 2 1059 1039
0 3030 7 1 2 1060 1045
0 3031 5 1 1 1296
0 3032 5 1 1 1298
0 3033 5 1 1 1300
0 3034 5 1 1 1302
0 3035 9 2 1 1048
0 3038 9 2 1 1049
0 3041 5 10 1 1089
0 3052 5 10 1 1101
0 3063 5 4 1 1108
0 3068 5 2 1 1113
0 3071 7 1 2 98 1109
0 3072 7 1 2 95 1110
0 3073 7 1 2 99 1111
0 3074 7 1 2 96 1112
0 3075 5 10 1 1121
0 3086 5 10 1 1132
0 3097 5 10 1 1165
0 3108 5 10 1 1172
0 3119 5 10 1 1180
0 3130 5 10 1 1188
0 3141 5 1 1 1313
0 3142 5 1 1 1316
0 3143 5 1 1 1318
0 3144 5 1 1 1320
0 3145 5 1 1 1322
0 3146 5 1 1 1324
0 3147 5 10 1 1194
0 3158 5 10 1 1201
0 3169 5 10 1 1207
0 3180 5 10 1 1215
0 3191 9 2 1 1225
0 3194 5 1 1 1305
0 3195 5 1 1 1307
0 3196 5 1 1 1309
0 3197 5 1 1 1311
0 3198 5 1 1 1326
0 3199 5 1 1 1329
0 3200 9 2 1 924
0 3203 5 1 1 1331
3 3357 9 0 1 1392
3 3358 9 0 1 1394
3 3359 9 0 1 1395
3 3360 9 0 1 1397
0 3401 7 1 3 462 655 2824
0 3402 7 1 3 473 656 2826
0 3403 7 1 3 427 657 2828
0 3404 7 1 3 440 658 2830
0 3405 7 1 2 644 2823
0 3406 7 1 2 645 2825
0 3407 7 1 2 646 2827
0 3408 7 1 2 647 2829
0 3409 7 1 3 394 659 2840
0 3410 7 1 3 405 660 2842
0 3411 7 1 3 416 661 2844
0 3412 7 1 3 379 662 2846
0 3413 7 1 2 648 2839
0 3414 7 1 2 649 2841
0 3415 7 1 2 650 2843
0 3416 7 1 2 651 2845
0 3444 7 1 2 788 2902
0 3445 7 1 3 484 789 2904
0 3446 7 1 3 495 790 2906
0 3447 7 1 2 1072 2901
0 3448 7 1 2 1073 2903
0 3449 7 1 2 1074 2905
0 3450 7 1 3 508 663 2914
0 3451 7 1 3 528 664 2916
0 3452 7 1 3 539 665 2918
0 3453 7 1 2 652 2913
0 3454 7 1 2 653 2915
0 3455 7 1 2 654 2917
0 3456 7 2 2 2920 2350
0 3459 7 1 3 395 791 2927
0 3460 7 1 3 406 792 2929
0 3461 7 1 3 417 793 2931
0 3462 7 1 3 380 794 2933
0 3463 7 1 2 1075 2926
0 3464 7 1 2 1076 2928
0 3465 7 1 2 1077 2930
0 3466 7 1 2 1078 2932
0 3481 7 1 3 509 799 2974
0 3482 5 1 1 2980
0 3483 7 1 3 529 800 2976
0 3484 7 1 3 540 801 2978
0 3485 7 1 2 780 2973
0 3486 7 1 2 781 2975
0 3487 7 1 2 782 2977
0 3488 7 1 2 802 2988
0 3489 7 1 3 485 803 2990
0 3490 7 1 3 496 804 2992
0 3491 7 1 2 783 2987
0 3492 7 1 2 784 2989
0 3493 7 1 2 785 2991
0 3502 7 1 2 805 2999
0 3503 7 1 2 806 3006
0 3504 7 1 3 463 795 3016
0 3505 7 1 3 474 796 3018
0 3506 7 1 3 428 797 3020
0 3507 7 1 3 441 798 3022
0 3508 7 1 2 1079 3015
0 3509 7 1 2 1081 3017
0 3510 7 1 2 1082 3019
0 3511 7 1 2 1083 3021
0 3512 6 1 2 1299 3031
0 3513 6 1 2 1297 3032
0 3514 6 1 2 1304 3033
0 3515 6 1 2 1301 3034
0 3558 6 1 2 1317 3141
0 3559 6 1 2 1314 3142
0 3560 6 1 2 1321 3143
0 3561 6 1 2 1319 3144
0 3562 6 1 2 1325 3145
0 3563 6 1 2 1323 3146
3 3604 9 0 1 1741
0 3605 6 1 2 1308 3194
0 3606 6 1 2 1306 3195
0 3607 6 1 2 1312 3196
0 3608 6 1 2 1310 3197
0 3609 6 1 2 1330 3198
0 3610 6 1 2 1328 3199
3 3613 5 0 1 1742
0 3614 7 1 2 1528 1536
0 3615 7 1 2 931 1537
0 3616 7 1 3 201 1338 698
0 3617 7 1 3 204 1340 699
0 3618 7 1 3 198 1341 700
0 3619 7 1 3 195 1342 701
0 3620 7 1 3 192 1343 702
0 3621 7 1 3 183 1366 721
0 3622 7 1 3 189 1367 722
0 3623 7 1 3 156 1368 723
0 3624 7 1 3 150 1369 724
0 3625 7 1 2 1529 1538
0 3626 7 1 2 932 1539
0 3627 7 1 3 202 1403 753
0 3628 7 1 3 205 1404 754
0 3629 7 1 3 199 1405 755
0 3630 7 1 3 196 1406 756
0 3631 7 1 3 193 1407 757
0 3632 7 1 3 184 1435 775
0 3633 7 1 3 190 1437 776
0 3634 7 1 3 157 1438 777
0 3635 7 1 3 151 1439 778
0 3636 7 1 2 1530 1540
0 3637 7 1 2 933 1541
0 3638 7 1 3 110 1619 1133
0 3639 7 1 2 1531 1543
0 3640 7 1 2 934 1544
0 3641 7 1 3 12 1457 849
0 3642 7 1 3 111 1582 1102
0 3643 7 1 3 47 1584 1103
0 3644 7 1 3 101 1585 1105
0 3645 7 1 3 92 1586 1106
0 3646 7 1 3 44 1587 1107
0 3647 7 1 3 77 1458 850
0 3648 7 1 3 74 1459 851
0 3649 7 1 3 68 1460 852
0 3650 7 1 3 15 1461 853
0 3651 7 1 3 48 1620 1134
0 3652 7 1 3 102 1622 1135
0 3653 7 1 3 93 1623 1136
0 3654 7 1 3 45 1625 1158
0 3655 7 1 3 78 1481 871
0 3656 7 1 3 75 1483 872
0 3657 7 1 3 69 1484 873
0 3658 7 1 3 16 1485 874
0 3659 7 1 3 120 1674 1189
0 3660 7 1 3 13 1486 875
0 3661 7 1 3 118 1649 1174
0 3662 7 1 3 177 1370 725
0 3663 7 1 3 178 1440 779
0 3664 3 1 2 2831 3401
0 3665 3 1 2 2832 3402
0 3666 3 1 2 2833 3403
0 3667 3 1 2 2834 3404
0 3668 3 1 3 2835 3405 464
0 3669 3 1 3 2836 3406 475
0 3670 3 1 3 2837 3407 429
0 3671 3 1 3 2838 3408 442
0 3672 3 1 2 2847 3409
0 3673 3 1 2 2848 3410
0 3674 3 1 2 2849 3411
0 3675 3 1 2 2850 3412
0 3676 3 1 3 2851 3413 396
0 3677 3 1 3 2852 3414 407
0 3678 3 1 3 2853 3415 418
0 3679 3 1 3 2854 3416 381
0 3680 7 1 2 291 1508
0 3681 7 1 2 287 1509
0 3682 7 1 2 279 1511
0 3683 7 1 2 271 1512
0 3684 7 1 2 263 1514
0 3685 7 1 2 240 1515
0 3686 7 1 2 232 1517
0 3687 7 1 2 224 1518
0 3688 7 1 2 216 1520
0 3689 7 1 2 208 1521
0 3691 5 8 1 1546
0 3700 3 1 2 2907 3444
0 3701 3 1 2 2908 3445
0 3702 3 1 2 2909 3446
0 3703 3 1 3 2911 3448 486
0 3704 3 1 3 2912 3449 497
0 3705 3 2 2 2910 3447
0 3708 3 1 2 2919 3450
0 3709 3 1 2 2921 3451
0 3710 3 1 2 2922 3452
0 3711 3 1 3 2923 3453 510
0 3712 3 1 3 2924 3454 530
0 3713 3 1 3 2925 3455 541
0 3715 3 1 2 2934 3459
0 3716 3 1 2 2935 3460
0 3717 3 1 2 2936 3461
0 3718 3 1 2 2937 3462
0 3719 3 1 3 2938 3463 397
0 3720 3 1 3 2939 3464 408
0 3721 3 1 3 2940 3465 419
0 3722 3 1 3 2941 3466 382
0 3723 7 1 2 371 1547
0 3724 7 1 2 365 1549
0 3725 7 1 2 357 1550
0 3726 7 1 2 347 1552
0 3727 7 1 2 330 1555
0 3728 7 1 2 322 1556
0 3729 7 1 2 314 1558
0 3730 7 1 2 306 1559
0 3731 7 1 2 298 1561
0 3732 3 5 2 1553 2958
0 3738 7 1 2 85 1562
0 3739 7 1 2 87 1564
0 3740 7 1 2 35 1565
0 3741 7 1 2 36 1567
0 3742 3 1 2 2979 3481
0 3743 3 1 2 2981 3483
0 3744 3 1 2 2982 3484
0 3745 3 1 3 2983 3485 511
0 3746 3 1 3 2985 3486 531
0 3747 3 1 3 2986 3487 542
0 3748 3 1 2 2993 3488
0 3749 3 1 2 2994 3489
0 3750 3 1 2 2995 3490
0 3751 3 1 3 2997 3492 487
0 3752 3 1 3 2998 3493 498
0 3753 5 1 1 1568
0 3754 5 1 1 1570
0 3755 5 1 1 1572
0 3756 5 1 1 1575
0 3757 3 1 2 3013 3502
0 3758 7 1 3 830 449 1571
0 3759 3 1 2 3014 3503
0 3760 7 1 3 831 450 1576
0 3761 7 1 2 1070 1569
0 3762 7 1 2 1071 1574
0 3763 3 1 2 3023 3504
0 3764 3 1 2 3024 3505
0 3765 3 1 2 3025 3506
0 3766 3 1 2 3026 3507
0 3767 3 1 3 3027 3508 465
0 3768 3 1 3 3028 3509 476
0 3769 3 1 3 3029 3510 430
0 3770 3 1 3 3030 3511 443
0 3771 6 3 2 3512 3513
0 3775 6 3 2 3514 3515
0 3779 5 1 1 1577
0 3780 5 1 1 1579
0 3781 7 1 3 117 1650 1175
0 3782 7 1 3 126 1652 1176
0 3783 7 1 3 127 1653 1177
0 3784 7 1 3 128 1655 1178
0 3785 7 1 3 131 1676 1190
0 3786 7 1 3 129 1677 1191
0 3787 7 1 3 119 1678 1192
0 3788 7 1 3 130 1679 1193
0 3789 6 3 2 3558 3559
0 3793 6 3 2 3560 3561
0 3797 6 2 2 3562 3563
0 3800 7 1 3 122 1696 1202
0 3801 7 1 3 113 1698 1203
0 3802 7 1 3 53 1699 1204
0 3803 7 1 3 114 1700 1205
0 3804 7 1 3 115 1701 1206
0 3805 7 1 3 52 1718 1217
0 3806 7 1 3 112 1719 1218
0 3807 7 1 3 116 1720 1220
0 3808 7 1 3 121 1722 1221
0 3809 7 1 3 125 1723 1222
0 3810 6 2 2 3607 3608
0 3813 6 2 2 3605 3606
0 3816 7 2 2 3482 2984
0 3819 3 2 2 2996 3491
0 3822 5 1 1 1744
0 3823 6 1 2 1745 3203
0 3824 6 2 2 3609 3610
0 3827 5 1 1 1746
0 3828 3 1 2 3739 2970
0 3829 3 1 2 3740 2971
0 3830 3 1 2 3741 2972
0 3831 3 1 2 3738 2969
0 3834 5 1 1 3664
0 3835 5 1 1 3665
0 3836 5 1 1 3666
0 3837 5 1 1 3667
0 3838 5 1 1 3672
0 3839 5 1 1 3673
0 3840 5 1 1 3674
0 3841 5 1 1 3675
0 3842 3 6 2 3681 2868
0 3849 3 5 2 3682 2869
0 3855 3 5 2 3683 2870
0 3861 3 5 2 3684 2871
0 3867 3 5 2 3685 2872
0 3873 3 7 2 3686 2873
0 3881 3 5 2 3687 2874
0 3887 3 5 2 3688 2875
0 3893 3 5 2 3689 2876
0 3908 5 1 1 3701
0 3909 5 1 1 3702
0 3911 5 2 1 3700
0 3914 5 1 1 3708
0 3915 5 1 1 3709
0 3916 5 1 1 3710
0 3917 5 1 1 3715
0 3918 5 1 1 3716
0 3919 5 1 1 3717
0 3920 5 1 1 3718
0 3921 3 5 2 3724 2955
0 3927 3 5 2 3725 2956
0 3933 3 5 2 3726 2957
0 3942 3 5 2 3727 2959
0 3948 3 7 2 3728 2960
0 3956 3 5 2 3729 2961
0 3962 3 5 2 3730 2962
0 3968 3 6 2 3731 2963
0 3975 5 1 1 3742
0 3976 5 1 1 3743
0 3977 5 1 1 3744
0 3978 5 1 1 3749
0 3979 5 1 1 3750
0 3980 7 1 3 451 807 3754
0 3981 7 1 3 452 808 3756
0 3982 7 1 2 786 3753
0 3983 7 1 2 787 3755
0 3984 5 2 1 3757
0 3987 5 1 1 3759
0 3988 5 1 1 3763
0 3989 5 1 1 3764
0 3990 5 1 1 3765
0 3991 5 1 1 3766
0 3998 7 1 3 1747 1680 1686
0 4008 3 2 2 3723 2954
0 4011 3 2 2 3680 2867
0 4021 5 2 1 3748
0 4024 6 1 2 1332 3822
0 4027 5 1 1 1757
0 4031 7 1 2 3828 993
0 4032 7 1 3 24 1532 1748
0 4033 7 1 3 25 935 1749
0 4034 7 1 3 26 1533 1750
0 4035 7 1 3 81 936 1751
0 4036 7 1 2 3829 994
0 4037 7 1 3 79 1534 1752
0 4038 7 1 3 23 937 1753
0 4039 7 1 3 82 1535 1754
0 4040 7 1 3 80 938 1756
0 4041 7 1 2 3830 995
0 4042 7 1 2 3831 996
0 4067 7 2 2 1760 521
0 4080 7 3 2 522 1762
0 4088 7 2 2 3834 3668
0 4091 7 2 2 3835 3669
0 4094 7 2 2 3836 3670
0 4097 7 2 2 3837 3671
0 4100 7 2 2 3838 3676
0 4103 7 2 2 3839 3677
0 4106 7 2 2 3840 3678
0 4109 7 2 2 3841 3679
0 4144 7 2 2 3908 3703
0 4147 7 2 2 3909 3704
0 4150 9 2 1 1759
0 4153 7 2 2 3914 3711
0 4156 7 2 2 3915 3712
0 4159 7 2 2 3916 3713
0 4183 3 1 2 3758 3980
0 4184 3 1 2 3760 3981
0 4185 3 1 3 3761 3982 453
0 4186 3 1 3 3762 3983 454
0 4188 5 2 1 1766
0 4191 5 2 1 1770
0 4196 7 1 3 1771 1767 1578
0 4197 7 1 3 3987 1681 1687
0 4198 7 1 2 3920 3722
0 4199 5 1 1 1787
0 4200 5 2 1 1773
0 4203 5 2 1 1776
0 4206 9 2 1 1780
0 4209 9 2 1 1781
0 4212 9 2 1 1763
0 4215 9 2 1 1764
0 4219 9 2 1 1765
0 4223 5 1 1 1782
0 4224 5 1 1 1784
0 4225 7 2 2 3918 3720
0 4228 7 2 2 3919 3721
0 4231 7 2 2 3991 3770
0 4234 7 2 2 3917 3719
0 4237 7 2 2 3989 3768
0 4240 7 2 2 3990 3769
0 4243 7 2 2 3988 3767
0 4246 7 2 2 3976 3746
0 4249 7 2 2 3977 3747
0 4252 7 2 2 3975 3745
0 4255 7 2 2 3978 3751
0 4258 7 2 2 3979 3752
0 4263 5 1 1 1789
0 4264 6 2 2 4024 3823
0 4267 5 1 1 1791
0 4268 7 1 2 455 1850
0 4269 5 1 1 1858
0 4270 5 1 1 1925
0 4271 7 1 2 1852 456
3 4272 5 0 1 4031
0 4273 3 1 4 4032 4033 3614 3615
0 4274 3 1 4 4034 4035 3625 3626
3 4275 5 0 1 4036
0 4276 3 1 4 4037 4038 3636 3637
0 4277 3 1 4 4039 4040 3639 3640
3 4278 5 0 1 4041
3 4279 5 0 1 4042
0 4280 7 3 2 1843 466
0 4284 7 5 2 1835 477
0 4290 7 6 2 431 1825
0 4297 7 1 2 1818 444
0 4298 7 2 2 1812 398
0 4301 7 3 2 1806 409
0 4305 7 4 2 1801 420
0 4310 7 5 2 1794 383
0 4316 7 3 2 467 1844
0 4320 7 4 2 478 1837
0 4325 7 5 2 432 1826
0 4331 7 1 2 445 1819
0 4332 7 3 2 399 1813
0 4336 7 5 2 410 1808
0 4342 7 6 2 421 1802
0 4349 7 7 2 384 1795
0 4357 5 6 1 1916
0 4364 5 10 1 1909
0 4375 9 3 1 1910
0 4379 7 5 2 1901 488
0 4385 7 6 2 499 1891
0 4392 7 1 2 1883 512
0 4396 7 3 2 1876 532
0 4400 7 4 2 1868 543
0 4405 5 6 1 1861
0 4412 9 5 1 1862
0 4418 5 6 1 1918
0 4425 5 10 1 1912
0 4436 9 3 1 1913
0 4440 7 4 2 489 1903
0 4445 7 5 2 500 1892
0 4451 7 1 2 513 1885
0 4456 7 5 2 533 1877
0 4462 7 6 2 544 1870
0 4469 9 7 1 1864
0 4477 5 6 1 1865
0 4512 9 2 1 1919
0 4515 5 1 1 4183
0 4516 5 1 1 4184
0 4521 5 1 1 1928
0 4523 5 1 1 1931
0 4524 5 3 1 4198
0 4532 5 3 1 1927
0 4547 7 1 3 1859 1724 1730
0 4548 9 2 1 1853
0 4551 9 2 1 1846
0 4554 9 2 1 1838
0 4557 9 2 1 1828
0 4560 9 2 1 1820
0 4563 9 2 1 1815
0 4566 9 2 1 1809
0 4569 9 2 1 1803
0 4572 9 2 1 1796
0 4575 4 2 2 433 1829
0 4578 9 2 1 1855
0 4581 9 2 1 1847
0 4584 9 2 1 1840
0 4587 9 2 1 1822
0 4590 9 2 1 1816
0 4593 9 2 1 1810
0 4596 9 2 1 1804
0 4599 9 2 1 1831
0 4602 9 2 1 1797
0 4605 4 2 2 434 1832
0 4608 4 2 2 385 1798
0 4611 9 2 1 1904
0 4614 9 2 1 1894
0 4617 9 2 1 1886
0 4621 9 2 1 1879
0 4624 9 2 1 1871
0 4627 4 2 2 501 1895
0 4630 9 2 1 1906
0 4633 9 2 1 1888
0 4637 9 2 1 1880
0 4640 9 2 1 1873
0 4643 9 2 1 1897
0 4646 4 2 2 502 1898
0 4649 9 2 1 1874
0 4652 9 2 1 1882
0 4655 9 2 1 1867
0 4658 9 2 1 1889
0 4662 9 2 1 1907
0 4665 9 2 1 1900
0 4668 9 2 1 1921
0 4671 9 2 1 1915
0 4674 9 2 1 1834
0 4677 9 2 1 1823
0 4680 9 2 1 1849
0 4683 9 2 1 1841
0 4686 9 2 1 1856
0 4689 9 2 1 1805
0 4692 9 2 1 1799
0 4695 9 2 1 1817
0 4698 9 2 1 1811
0 4701 6 1 2 1786 4223
0 4702 6 1 2 1783 4224
0 4720 5 1 1 1934
0 4721 6 1 2 1936 4263
0 4724 5 1 1 1971
0 4725 5 1 1 1969
0 4726 5 1 1 1980
0 4727 5 1 1 1978
0 4728 5 1 1 1976
0 4729 5 1 1 1954
0 4730 5 1 1 1951
0 4731 5 1 1 1948
0 4732 5 1 1 1945
0 4733 5 1 1 1966
0 4734 5 1 1 1963
0 4735 5 1 1 1960
0 4736 5 1 1 1957
3 4737 7 0 2 4273 1523
3 4738 7 0 2 4274 1524
3 4739 7 0 2 4276 1526
3 4740 7 0 2 4277 1527
0 4741 7 1 3 1974 1163 1159
0 4855 5 1 1 1994
0 4856 6 1 2 1995 2712
0 4908 6 1 2 1996 2718
0 4909 5 1 1 1997
0 4939 7 2 2 4515 4185
0 4942 7 1 2 4516 4186
0 4947 5 1 1 1998
0 4953 7 1 3 1982 1772 3779
0 4954 7 1 3 1768 1984 3780
0 4955 7 1 3 1985 1983 1581
0 4956 7 1 3 1967 1656 1664
0 4957 7 1 3 1964 1658 1665
0 4958 7 1 3 1961 1659 1666
0 4959 7 1 3 1958 1661 1667
0 4960 7 1 3 1981 1682 1688
0 4961 7 1 3 1979 1683 1689
0 4965 5 1 1 2000
0 4966 5 1 1 2002
0 4967 5 1 1 2004
0 4968 5 1 1 2006
0 4972 5 1 1 2014
0 4973 5 1 1 2016
0 4974 5 1 1 2018
0 4975 6 1 2 2019 4199
0 4976 5 1 1 1990
0 4977 5 1 1 1992
0 4978 7 1 3 1778 1774 1991
0 4979 7 1 3 1988 1986 1993
0 4980 7 1 3 1955 1702 1707
0 4981 7 1 3 1952 1703 1708
0 4982 7 1 3 1949 1704 1710
0 4983 7 1 3 1946 1705 1711
0 4984 7 1 3 1977 1725 1732
0 4985 7 1 3 1973 1726 1733
0 4986 7 1 3 1970 1728 1734
0 4987 7 1 3 1975 1729 1735
0 5049 6 2 2 4701 4702
0 5052 5 1 1 2008
0 5053 5 1 1 2010
0 5054 5 1 1 2012
0 5055 5 1 1 2020
0 5056 5 1 1 2022
0 5057 6 1 2 1790 4720
0 5058 5 1 1 2024
0 5059 6 1 2 2025 4267
0 5060 7 1 4 4724 4725 4269 4027
0 5061 7 1 4 4726 4727 3827 4728
0 5062 7 1 4 4729 4730 4731 4732
0 5063 7 1 4 4733 4734 4735 4736
0 5065 7 1 2 2090 2106
0 5066 7 1 3 2096 2091 2109
0 5067 7 1 2 2138 2156
0 5068 7 1 3 2146 2140 2159
0 5069 5 1 1 2200
0 5070 6 1 2 2201 2628
0 5071 5 1 1 2202
0 5072 6 1 2 2203 2629
0 5073 5 1 1 2204
0 5074 6 1 2 2205 2630
0 5075 5 1 1 2206
0 5076 6 1 2 2207 2631
0 5077 5 1 1 2208
0 5078 6 1 2 2209 2632
0 5079 5 1 1 2210
0 5080 6 1 2 2211 2633
0 5081 5 1 1 2212
0 5082 6 1 2 2213 2634
0 5083 5 1 1 2214
0 5084 6 1 2 2215 2635
0 5085 5 1 1 2216
0 5086 6 1 2 2217 2636
0 5087 5 1 1 2218
0 5088 6 1 2 2220 2638
0 5089 5 1 1 2221
0 5090 6 1 2 2222 2639
0 5091 5 1 1 2223
0 5092 6 1 2 2224 2640
0 5093 5 1 1 2225
0 5094 6 1 2 2226 2641
0 5095 5 1 1 2227
0 5096 6 1 2 2228 2642
0 5097 5 1 1 2229
0 5098 6 1 2 2230 2643
0 5099 5 1 1 2231
0 5100 6 1 2 2232 2644
0 5101 5 1 1 2233
0 5102 6 1 2 2234 2645
0 5103 5 1 1 2235
0 5104 6 1 2 2236 2646
0 5105 5 1 1 2237
0 5106 5 1 1 2242
0 5107 6 1 2 2243 2709
0 5108 5 1 1 2244
0 5109 6 1 2 2245 2710
0 5110 5 1 1 2246
0 5111 6 1 2 2247 2711
0 5112 6 1 2 1275 4855
0 5113 5 1 1 2248
0 5114 6 1 2 2249 2713
0 5115 5 1 1 2250
0 5116 6 1 2 2251 2714
0 5117 7 1 2 2097 2110
0 5118 7 1 2 2098 2111
0 5119 7 1 2 56 2127
0 5120 5 1 1 2252
0 5121 6 1 2 2254 2716
0 5122 5 1 1 2255
0 5123 6 1 2 2256 2717
0 5124 5 1 1 2257
0 5125 6 1 2 1288 4909
0 5126 6 1 2 2258 2719
0 5127 5 1 1 2259
0 5128 6 1 2 2260 2720
0 5129 5 1 1 2261
0 5130 6 1 2 2262 2721
0 5131 5 1 1 2263
0 5132 7 1 2 2147 2160
0 5133 7 1 2 2148 2161
0 5135 5 1 1 2266
0 5136 5 1 1 2268
0 5137 6 1 2 2270 4521
0 5138 5 1 1 2271
0 5139 5 1 1 2272
0 5140 6 1 2 2273 4947
0 5141 5 1 1 2282
0 5142 5 1 1 2284
0 5143 5 1 1 2286
0 5144 5 1 1 2288
0 5145 6 1 2 2290 4523
0 5146 5 1 1 2291
0 5147 4 1 2 4953 4196
0 5148 4 1 2 4954 4955
0 5150 5 2 1 2194
0 5153 6 1 2 2003 4965
0 5154 6 1 2 2001 4966
0 5155 6 1 2 2007 4967
0 5156 6 1 2 2005 4968
0 5157 5 2 1 2197
0 5160 6 1 2 2017 4972
0 5161 6 1 2 2015 4973
0 5162 6 1 2 1788 4974
0 5163 7 1 3 1987 1779 4976
0 5164 7 1 3 1775 1989 4977
0 5165 7 1 3 4942 1706 1712
0 5166 5 2 1 2192
0 5169 9 2 1 2034
0 5172 5 1 1 2238
0 5173 9 2 1 2064
0 5176 5 1 1 2240
0 5177 9 2 1 2083
0 5180 9 2 1 2128
0 5183 9 2 1 2092
0 5186 9 2 1 2093
0 5189 9 2 1 2099
0 5192 9 2 1 2100
0 5195 9 2 1 2114
0 5198 5 1 1 2264
0 5199 9 2 1 2141
0 5202 9 2 1 2149
0 5205 9 2 1 2163
0 5208 9 2 1 2143
0 5211 9 2 1 2150
0 5214 9 2 1 2186
0 5217 9 2 1 2179
0 5220 9 2 1 2187
0 5223 5 1 1 2274
0 5224 5 1 1 2276
0 5225 5 1 1 2278
0 5226 5 1 1 2280
0 5227 5 1 1 2292
0 5228 5 1 1 2294
0 5229 5 1 1 2296
0 5230 5 1 1 2298
0 5232 6 1 2 2011 5052
0 5233 6 1 2 2009 5053
0 5234 6 1 2 2023 5055
0 5235 6 1 2 2021 5056
0 5236 6 2 2 4721 5057
0 5239 6 1 2 1792 5058
3 5240 7 0 3 5060 5061 4270
0 5241 5 1 1 2300
0 5242 6 1 2 1227 5069
0 5243 6 1 2 1229 5071
0 5244 6 1 2 1231 5073
0 5245 6 1 2 1233 5075
0 5246 6 1 2 1236 5077
0 5247 6 1 2 1238 5079
0 5248 6 1 2 1240 5081
0 5249 6 1 2 1242 5083
0 5250 6 1 2 1244 5085
0 5252 6 1 2 1249 5089
0 5253 6 1 2 1251 5091
0 5254 6 1 2 1253 5093
0 5255 6 1 2 1255 5095
0 5256 6 1 2 1257 5097
0 5257 6 1 2 1260 5099
0 5258 6 1 2 1262 5101
0 5259 6 1 2 1264 5103
0 5260 6 1 2 1266 5105
0 5261 6 1 2 1268 5106
0 5262 6 1 2 1270 5108
0 5263 6 1 2 1273 5110
0 5264 6 9 2 5112 4856
0 5274 6 1 2 1277 5113
0 5275 6 1 2 1279 5115
0 5282 6 1 2 1284 5122
0 5283 6 1 2 1286 5124
0 5284 6 13 2 4908 5125
0 5298 6 1 2 1290 5127
0 5299 6 1 2 1293 5129
0 5300 6 1 2 1295 5131
0 5303 6 1 2 2269 5135
0 5304 6 1 2 2267 5136
0 5305 6 1 2 1930 5138
0 5306 6 1 2 1999 5139
0 5307 6 1 2 2285 5141
0 5308 6 1 2 2283 5142
0 5309 6 1 2 2289 5143
0 5310 6 1 2 2287 5144
0 5311 6 1 2 1933 5146
0 5312 5 1 1 2302
0 5315 6 3 2 5153 5154
0 5319 6 2 2 5155 5156
0 5324 6 3 2 5160 5161
0 5328 6 2 2 5162 4975
0 5331 4 1 2 5163 4978
0 5332 4 1 2 5164 4979
0 5346 3 2 2 2133 5119
0 5363 6 1 2 2277 5223
0 5364 6 1 2 2275 5224
0 5365 6 1 2 2281 5225
0 5366 6 1 2 2279 5226
0 5367 6 1 2 2295 5227
0 5368 6 1 2 2293 5228
0 5369 6 1 2 2299 5229
0 5370 6 1 2 2297 5230
0 5371 6 2 2 5148 5147
0 5374 9 2 1 2301
0 5377 6 2 2 5232 5233
0 5382 6 2 2 5234 5235
0 5385 6 2 2 5239 5059
3 5388 7 0 3 5062 5063 5241
0 5389 6 6 2 5242 5070
0 5396 6 10 2 5243 5072
0 5407 6 10 2 5244 5074
0 5418 6 5 2 5245 5076
0 5424 6 6 2 5246 5078
0 5431 6 9 2 5247 5080
0 5441 6 10 2 5248 5082
0 5452 6 9 2 5249 5084
0 5462 6 6 2 5250 5086
0 5469 5 1 1 2311
0 5470 6 6 2 5088 5252
0 5477 6 10 2 5090 5253
0 5488 6 9 2 5092 5254
0 5498 6 7 2 5094 5255
0 5506 6 13 2 5096 5256
0 5520 6 15 2 5098 5257
0 5536 6 12 2 5100 5258
0 5549 6 5 2 5102 5259
0 5555 6 6 2 5104 5260
0 5562 6 10 2 5261 5107
0 5573 6 5 2 5262 5109
0 5579 6 6 2 5263 5111
0 5595 6 10 2 5274 5114
0 5606 6 9 2 5275 5116
0 5616 6 1 2 2317 2715
0 5617 5 1 1 2318
0 5618 5 1 1 2319
0 5619 5 1 1 2321
0 5620 5 1 1 2323
0 5621 5 1 1 2325
0 5622 5 1 1 2327
0 5624 6 9 2 5121 5282
0 5634 6 7 2 5123 5283
0 5655 6 15 2 5126 5298
0 5671 6 12 2 5128 5299
0 5684 6 5 2 5130 5300
0 5690 5 1 1 2331
0 5691 5 1 1 2337
0 5692 6 3 2 5303 5304
0 5696 6 3 2 5137 5305
0 5700 6 2 2 5306 5140
0 5703 6 3 2 5307 5308
0 5707 6 3 2 5309 5310
0 5711 6 2 2 5145 5311
0 5726 7 1 2 2308 2193
0 5727 5 1 1 2313
0 5728 5 1 1 2315
0 5730 5 1 1 2329
0 5731 5 1 1 2333
0 5732 5 1 1 2335
0 5733 5 1 1 2339
0 5734 5 1 1 2341
0 5735 5 1 1 2343
0 5736 6 2 2 5365 5366
0 5739 6 2 2 5363 5364
0 5742 6 2 2 5369 5370
0 5745 6 2 2 5367 5368
0 5755 5 1 1 2345
0 5756 6 2 2 5332 5331
0 5954 7 1 2 2347 2120
0 5955 6 1 2 1282 5617
0 5956 5 1 1 2381
0 6005 7 1 2 2358 2168
0 6006 7 1 2 2359 2169
0 6023 5 1 1 2383
0 6024 6 1 2 2384 5312
0 6025 5 2 1 2371
0 6028 5 2 1 2376
0 6031 9 2 1 2374
0 6034 9 2 1 2375
0 6037 9 2 1 2379
0 6040 9 2 1 2380
0 6044 5 1 1 2392
0 6045 3 2 2 2310 5726
0 6048 9 2 1 2348
0 6051 9 2 1 2360
0 6054 9 2 1 2361
0 6065 5 1 1 2385
0 6066 6 1 2 2386 5054
0 6067 5 1 1 2388
0 6068 5 1 1 2390
0 6069 6 1 2 2391 5755
0 6071 7 1 2 2465 2055
0 6072 7 1 3 2471 2466 2058
0 6073 7 1 4 2481 2467 2065 2472
0 6074 7 1 4 2549 2094 2115 2101
0 6075 7 1 2 2394 2026
0 6076 7 1 3 2400 2395 2029
0 6077 7 1 4 2410 2396 2035 2401
0 6078 7 1 4 2654 2144 2164 2151
0 6079 5 1 1 2420
0 6080 7 2 4 2402 2421 2411 2397
0 6083 7 1 2 2403 2030
0 6084 7 1 3 2412 2036 2404
0 6085 7 1 3 2422 2413 2405
0 6086 7 1 2 2406 2031
0 6087 7 1 3 2037 2414 2407
0 6088 7 1 2 2415 2038
0 6089 7 1 2 2423 2416
0 6090 7 1 2 2417 2039
0 6091 7 2 5 2431 2459 2440 2425 2450
0 6094 7 1 2 2426 2040
0 6095 7 1 3 2432 2427 2042
0 6096 7 1 4 2441 2428 2045 2433
0 6097 7 1 5 2451 2442 2429 2049 2434
0 6098 7 1 2 2435 2043
0 6099 7 1 3 2443 2046 2436
0 6100 7 1 4 2452 2444 2050 2437
0 6101 7 1 5 6 2460 2445 2453 2438
0 6102 7 1 2 2047 2446
0 6103 7 1 3 2454 2447 2051
0 6104 7 1 4 7 2461 2448 2455
0 6105 7 1 2 2456 2052
0 6106 7 1 3 8 2462 2457
0 6107 7 1 2 9 2463
0 6108 7 2 4 2538 2482 2473 2468
0 6111 7 1 2 2474 2059
0 6112 7 1 3 2483 2066 2475
0 6113 7 1 3 2539 2484 2476
0 6114 7 1 2 2477 2062
0 6115 7 1 3 2485 2067 2478
0 6116 7 1 2 2486 2068
0 6117 7 2 5 2543 2525 2510 2497 2490
0 6120 7 1 2 2491 2069
0 6121 7 1 3 2498 2492 2072
0 6122 7 1 4 2511 2493 2077 2499
0 6123 7 1 5 2526 2512 2494 2084 2500
0 6124 7 1 2 2501 2073
0 6125 7 1 3 2513 2078 2502
0 6126 7 1 4 2528 2514 2085 2503
0 6127 7 1 4 2544 2515 2504 2529
0 6128 7 1 2 2505 2074
0 6129 7 1 3 2516 2079 2506
0 6130 7 1 4 2530 2517 2086 2507
0 6131 7 1 2 2518 2080
0 6132 7 1 3 2531 2519 2087
0 6133 7 1 3 2545 2520 2532
0 6134 7 1 2 2521 2081
0 6135 7 1 3 2533 2522 2088
0 6136 7 1 2 2534 2089
0 6137 7 1 2 2540 2487
0 6138 7 1 2 2546 2535
0 6139 5 1 1 2559
0 6140 7 2 4 2102 2560 2550 2095
0 6143 7 1 3 2551 2116 2103
0 6144 7 1 3 2561 2552 2104
0 6145 7 1 3 2117 2553 2105
0 6146 7 1 2 2554 2118
0 6147 7 1 2 2562 2555
0 6148 7 1 2 2556 2119
0 6149 7 2 5 2351 2129 2570 2564 2580
0 6152 7 1 2 2565 1937
0 6153 7 1 3 2352 2566 2121
0 6154 7 1 4 2571 2567 2123 2353
0 6155 7 1 5 2581 2572 2568 2134 2354
0 6156 7 1 3 2573 2124 2355
0 6157 7 1 4 2582 2574 2135 2356
0 6158 7 1 5 57 2130 2575 2583 2357
0 6159 7 1 2 2125 2576
0 6160 7 1 3 2648 2577 2136
0 6161 7 1 4 58 2131 2578 2649
0 6162 7 1 2 2650 2137
0 6163 7 1 3 59 2132 2651
0 6164 6 2 2 5616 5955
0 6168 7 2 4 2701 2655 2152 2145
0 6171 7 1 3 2656 2165 2153
0 6172 7 1 3 2702 2657 2154
0 6173 7 1 3 2658 2166 2155
0 6174 7 1 2 2659 2167
0 6175 7 2 5 2188 2688 2671 2362 2663
0 6178 7 1 2 2665 1940
0 6179 7 1 3 2363 2666 2170
0 6180 7 1 4 2672 2667 2173 2364
0 6181 7 1 5 2689 2673 2668 2180 2365
0 6182 7 1 3 2674 2174 2366
0 6183 7 1 4 2690 2676 2181 2367
0 6184 7 1 4 2189 2677 2368 2691
0 6185 7 1 3 2678 2175 2369
0 6186 7 1 4 2693 2679 2182 2370
0 6187 7 1 2 2680 2176
0 6188 7 1 3 2694 2682 2183
0 6189 7 1 3 2190 2683 2695
0 6190 7 1 2 2684 2177
0 6191 7 1 3 2696 2685 2184
0 6192 7 1 2 2697 2185
0 6193 7 1 2 2705 2660
0 6194 7 1 2 2191 2698
0 6197 5 2 1 2708
0 6200 5 2 1 2725
0 6203 5 2 1 2731
0 6206 5 2 1 2734
0 6209 9 2 1 2729
0 6212 9 2 1 2730
0 6215 9 2 1 2737
0 6218 9 2 1 2738
0 6221 6 1 2 2303 6023
0 6234 5 1 1 2748
0 6235 6 1 2 2749 6044
0 6238 9 2 1 2464
0 6241 9 2 1 2398
0 6244 9 2 1 2399
0 6247 9 2 1 2408
0 6250 9 2 1 2409
0 6253 9 2 1 2418
0 6256 9 2 1 2419
0 6259 9 2 1 2430
0 6262 9 2 1 2439
0 6265 9 2 1 2449
0 6268 9 2 1 2458
0 6271 9 2 1 2541
0 6274 9 2 1 2488
0 6277 9 2 1 2469
0 6280 9 2 1 2479
0 6283 9 2 1 2542
0 6286 9 2 1 2489
0 6289 9 2 1 2470
0 6292 9 2 1 2480
0 6295 9 2 1 2547
0 6298 9 2 1 2536
0 6301 9 2 1 2495
0 6304 9 2 1 2523
0 6307 9 2 1 2508
0 6310 9 2 1 2509
0 6313 9 2 1 2548
0 6316 9 2 1 2537
0 6319 9 2 1 2496
0 6322 9 2 1 2524
0 6325 9 2 1 2557
0 6328 9 2 1 2558
0 6331 9 2 1 2569
0 6335 9 2 1 2579
0 6338 9 2 1 2652
0 6341 9 2 1 2706
0 6344 9 2 1 2661
0 6347 9 2 1 2707
0 6350 9 2 1 2662
0 6353 9 2 1 2699
0 6356 9 2 1 2669
0 6359 9 2 1 2686
0 6364 9 2 1 2700
0 6367 9 2 1 2670
0 6370 9 2 1 2687
0 6373 5 1 1 2740
0 6374 5 1 1 2742
0 6375 5 1 1 2744
0 6376 5 1 1 2746
0 6377 6 1 2 2013 6065
0 6378 6 1 2 2346 6068
0 6382 3 1 4 4268 6071 6072 6073
0 6386 3 1 4 1922 5065 5066 6074
0 6388 3 1 4 4271 6075 6076 6077
0 6392 3 1 4 1924 5067 5068 6078
0 6397 3 2 5 4297 6094 6095 6096 6097
0 6411 3 2 2 2063 6116
0 6415 3 3 5 4331 6120 6121 6122 6123
0 6419 3 2 2 2082 6136
0 6427 3 2 5 4392 6152 6153 6154 6155
0 6434 5 1 1 2766
0 6437 3 2 2 2162 6174
0 6441 3 3 5 4451 6178 6179 6180 6181
0 6445 3 2 2 2178 6192
0 6448 5 1 1 2769
0 6449 5 1 1 2771
0 6466 6 2 2 6221 6024
0 6469 5 1 1 2755
0 6470 5 1 1 2758
0 6471 5 1 1 2760
0 6472 5 1 1 2762
0 6473 7 1 3 2372 2195 2757
0 6474 7 1 3 2751 2304 2759
0 6475 7 1 3 2377 2198 2761
0 6476 7 1 3 2753 2306 2763
0 6477 6 1 2 2393 6234
0 6478 6 2 2 2764 133
0 6482 3 2 4 2027 6083 6084 6085
0 6486 4 2 3 2028 6086 6087
0 6490 3 2 3 2032 6088 6089
0 6494 4 2 2 2033 6090
0 6500 3 2 5 2041 6098 6099 6100 6101
0 6504 3 2 4 2044 6102 6103 6104
0 6508 3 2 3 2048 6105 6106
0 6512 3 2 2 2053 6107
0 6516 3 2 4 2056 6111 6112 6113
0 6526 4 2 3 2057 6114 6115
0 6536 3 2 4 2075 6131 6132 6133
0 6539 3 2 5 2070 6124 6125 6126 6127
0 6553 4 2 3 2076 6134 6135
0 6556 4 2 4 2071 6128 6129 6130
0 6566 3 2 4 2107 5117 6143 6144
0 6569 4 2 3 2108 5118 6145
0 6572 3 2 3 2112 6146 6147
0 6575 4 2 2 2113 6148
0 6580 3 2 5 1939 5954 6156 6157 6158
0 6584 3 2 4 2122 6159 6160 6161
0 6587 3 2 3 2126 6162 6163
0 6592 3 2 4 2157 5132 6171 6172
0 6599 4 2 3 2158 5133 6173
0 6606 3 2 4 2171 6187 6188 6189
0 6609 3 2 5 1942 6005 6182 6183 6184
0 6619 4 2 3 2172 6190 6191
0 6622 4 2 4 1943 6006 6185 6186
0 6630 6 1 2 2743 6373
0 6631 6 1 2 2741 6374
0 6632 6 1 2 2747 6375
0 6633 6 1 2 2745 6376
0 6634 6 2 2 6377 6066
0 6637 6 2 2 6069 6378
0 6640 5 1 1 2787
3 6641 7 0 2 2777 2781
3 6643 7 0 2 2783 2785
3 6646 7 0 2 2789 2792
3 6648 7 0 2 2773 2775
0 6650 6 1 2 2811 2637
0 6651 5 1 1 2813
0 6653 5 1 1 2814
0 6655 5 1 1 2816
0 6657 5 1 1 2818
0 6659 5 1 1 2820
0 6660 6 1 2 2822 5087
0 6661 5 1 1 2856
0 6662 6 1 2 2857 5469
0 6663 5 1 1 2858
0 6664 7 1 2 2776 10
0 6666 5 1 1 2859
0 6668 5 1 1 2862
0 6670 5 1 1 2864
0 6672 5 1 1 2866
0 6675 5 1 1 2782
0 6680 5 1 1 2886
0 6681 5 1 1 2895
0 6682 5 1 1 2947
0 6683 5 1 1 2950
0 6689 6 1 2 3004 5120
0 6690 5 1 1 3005
0 6691 6 1 2 3008 5622
0 6692 5 1 1 3009
0 6693 7 1 2 2786 60
0 6695 5 1 1 3011
0 6698 5 1 1 3036
0 6699 6 1 2 3039 5956
0 6700 5 1 1 3040
0 6703 5 1 1 2793
0 6708 5 1 1 2803
0 6709 5 1 1 2805
0 6710 5 1 1 2807
0 6711 5 1 1 2809
0 6712 7 1 3 2726 2723 2804
0 6713 7 1 3 2796 2794 2806
0 6714 7 1 3 2735 2732 2808
0 6715 7 1 3 2800 2798 2810
3 6716 9 0 1 3089
0 6718 7 1 3 2788 1181 1690
0 6719 7 1 3 2305 2373 6469
0 6720 7 1 3 2196 2752 6470
0 6721 7 1 3 2307 2378 6471
0 6722 7 1 3 2199 2754 6472
0 6724 6 2 2 6477 6235
0 6739 5 1 1 2879
0 6740 5 1 1 2881
0 6741 5 1 1 2884
0 6744 5 1 1 2888
0 6745 5 1 1 2890
0 6746 5 1 1 2893
0 6751 5 1 1 2897
0 6752 5 1 1 2899
0 6753 5 1 1 2943
0 6754 5 1 1 2945
0 6755 5 1 1 3001
0 6760 5 1 1 2952
0 6761 5 1 1 2965
0 6762 5 1 1 2967
0 6772 5 1 1 3042
0 6773 5 1 1 3044
0 6776 5 1 1 3046
0 6777 5 1 1 3048
0 6782 5 1 1 3050
0 6783 5 1 1 3053
0 6784 5 1 1 3055
0 6785 5 1 1 3061
0 6790 5 1 1 3057
0 6791 5 1 1 3059
0 6792 6 2 2 6630 6631
0 6795 6 2 2 6632 6633
0 6801 7 1 2 2780 3069
0 6802 7 1 2 3079 2784
0 6803 7 1 2 3064 2774
0 6804 7 1 2 2791 3083
0 6805 5 1 1 3090
0 6806 6 1 2 1246 6651
0 6807 5 1 1 3093
0 6808 6 1 2 3094 6653
0 6809 5 1 1 3095
0 6810 6 1 2 3096 6655
0 6811 5 1 1 3098
0 6812 6 1 2 3099 6657
0 6813 5 1 1 3100
0 6814 6 1 2 3101 6659
0 6815 6 1 2 2219 6661
0 6816 6 1 2 2312 6663
0 6817 3 5 2 3065 6664
0 6823 5 1 1 3102
0 6824 6 1 2 3103 6666
0 6825 5 1 1 3104
0 6826 6 1 2 3105 6668
0 6827 5 1 1 3106
0 6828 6 1 2 3107 6670
0 6829 5 1 1 3109
0 6830 6 1 2 3110 6672
0 6831 5 2 1 3070
0 6834 5 1 1 3124
0 6835 6 1 2 3125 5618
0 6836 5 1 1 3126
0 6837 6 1 2 3127 5619
0 6838 5 1 1 3128
0 6839 6 1 2 3129 5620
0 6840 5 1 1 3131
0 6841 6 1 2 3132 5621
0 6842 6 1 2 2253 6690
0 6843 6 1 2 2328 6692
0 6844 3 5 2 3080 6693
0 6850 5 1 1 3133
0 6851 6 1 2 3134 6695
0 6852 5 1 1 3135
0 6853 6 1 2 3136 6434
0 6854 5 1 1 3137
0 6855 6 1 2 3138 6698
0 6856 6 1 2 2382 6700
0 6857 5 2 1 3084
0 6860 7 1 3 2795 2727 6708
0 6861 7 1 3 2724 2797 6709
0 6862 7 1 3 2799 2736 6710
0 6863 7 1 3 2733 2802 6711
0 6866 3 5 3 4197 6718 3785
0 6872 4 1 2 6719 6473
0 6873 4 1 2 6720 6474
0 6874 4 1 2 6721 6475
0 6875 4 1 2 6722 6476
0 6876 5 1 1 3161
3 6877 9 0 1 3163
0 6879 7 1 2 2765 3091
0 6880 7 1 2 3092 134
0 6881 3 2 2 3066 6137
0 6884 5 1 1 3111
0 6885 5 2 1 3067
0 6888 5 1 1 3113
0 6889 5 1 1 3115
0 6890 6 1 2 3116 5176
0 6891 3 2 2 3077 6138
0 6894 5 1 1 3117
0 6895 5 1 1 3120
0 6896 6 1 2 3121 5728
0 6897 5 2 1 3078
0 6900 5 1 1 3122
0 6901 3 2 2 3081 6193
0 6904 5 1 1 3139
0 6905 5 2 1 3082
0 6908 5 1 1 3148
0 6909 3 2 2 3087 6194
0 6912 5 1 1 3150
0 6913 5 1 1 3152
0 6914 5 1 1 3154
0 6915 6 1 2 3155 5734
0 6916 5 2 1 3088
0 6919 5 1 1 3156
0 6922 5 1 1 3159
0 6923 6 1 2 3160 6067
3 6924 3 0 2 6382 6801
3 6925 3 0 2 6386 6802
3 6926 3 0 2 6388 6803
3 6927 3 0 2 6392 6804
0 6930 5 1 1 3164
0 6932 6 2 2 6650 6806
0 6935 6 1 2 2815 6807
0 6936 6 1 2 2817 6809
0 6937 6 1 2 2819 6811
0 6938 6 1 2 2821 6813
0 6939 6 1 2 6660 6815
0 6940 6 1 2 6662 6816
0 6946 6 1 2 2860 6823
0 6947 6 1 2 2863 6825
0 6948 6 1 2 2865 6827
0 6949 6 1 2 2878 6829
0 6953 6 1 2 2320 6834
0 6954 6 1 2 2322 6836
0 6955 6 1 2 2324 6838
0 6956 6 1 2 2326 6840
0 6957 6 1 2 6689 6842
0 6958 6 1 2 6691 6843
0 6964 6 1 2 3012 6850
0 6965 6 1 2 2768 6852
0 6966 6 1 2 3037 6854
0 6967 6 2 2 6699 6856
0 6973 4 1 2 6860 6712
0 6974 4 1 2 6861 6713
0 6975 4 1 2 6862 6714
0 6976 4 1 2 6863 6715
0 6977 5 1 1 3165
0 6978 5 1 1 3167
0 6979 3 3 2 6879 6880
0 6987 6 1 2 2241 6889
0 6990 6 1 2 2316 6895
0 6999 6 1 2 2342 6914
0 7002 6 1 2 2389 6922
0 7003 6 2 2 6873 6872
0 7006 6 2 2 6875 6874
0 7011 7 1 3 3185 1371 1377
0 7012 7 1 3 3186 1441 1446
0 7013 7 1 3 3187 1463 1468
3 7015 5 0 1 3188
0 7016 7 1 3 3189 1487 1493
0 7018 6 1 2 6935 6808
0 7019 6 1 2 6936 6810
0 7020 6 1 2 6937 6812
0 7021 6 1 2 6938 6814
0 7022 5 1 1 6939
0 7023 5 4 1 3170
0 7028 6 2 2 6946 6824
0 7031 6 2 2 6947 6826
0 7034 6 2 2 6948 6828
0 7037 6 2 2 6949 6830
0 7040 7 1 2 3171 6079
0 7041 7 2 2 3175 6675
0 7044 6 1 2 6953 6835
0 7045 6 1 2 6954 6837
0 7046 6 1 2 6955 6839
0 7047 6 1 2 6956 6841
0 7048 5 1 1 6957
0 7049 5 4 1 3177
0 7054 6 2 2 6964 6851
0 7057 6 2 2 6965 6853
0 7060 6 2 2 6966 6855
0 7064 7 1 2 3178 6139
0 7065 7 2 2 3183 6703
0 7072 5 1 1 3190
0 7073 6 1 2 3192 5172
0 7074 5 1 1 3193
0 7075 6 1 2 3201 5727
0 7076 6 2 2 6890 6987
0 7079 5 1 1 3202
0 7080 6 2 2 6896 6990
0 7083 5 1 1 3205
0 7084 5 1 1 3207
0 7085 6 1 2 3208 5198
0 7086 5 1 1 3209
0 7087 6 1 2 3210 5731
0 7088 5 1 1 3211
0 7089 6 1 2 3212 6912
0 7090 6 2 2 6915 6999
0 7093 5 1 1 3213
0 7094 6 2 2 6974 6973
0 7097 6 2 2 6976 6975
0 7101 6 2 2 7002 6923
0 7105 5 1 1 3215
0 7110 5 1 1 3217
0 7114 7 1 3 3219 605 1160
0 7115 5 1 1 7019
0 7116 5 1 1 7021
0 7125 7 1 2 3172 7018
0 7126 7 1 2 3173 7020
0 7127 7 1 2 3174 7022
0 7130 5 1 1 7045
0 7131 5 1 1 7047
0 7139 7 1 2 3179 7044
0 7140 7 1 2 3181 7046
0 7141 7 1 2 3182 7048
0 7146 7 1 3 3216 1166 1668
0 7147 7 1 3 3218 1182 1691
0 7149 5 1 1 3222
0 7150 5 1 1 3224
0 7151 6 1 2 3225 6876
0 7152 6 1 2 2239 7072
0 7153 6 1 2 2314 7074
0 7158 6 1 2 2265 7084
0 7159 6 1 2 2334 7086
0 7160 6 1 2 3151 7088
0 7166 5 1 1 3236
0 7167 5 1 1 3234
0 7168 5 1 1 3232
0 7169 5 1 1 3230
0 7170 5 1 1 3248
0 7171 5 1 1 3246
0 7172 5 1 1 3244
0 7173 7 1 2 7115 3226
0 7174 7 1 2 7116 3227
0 7175 7 1 2 6940 3228
0 7176 7 1 2 2424 3229
0 7177 5 1 1 3238
0 7178 7 1 2 7130 3240
0 7179 7 1 2 7131 3241
0 7180 7 1 2 6958 3242
0 7181 7 1 2 2563 3243
0 7182 5 1 1 3250
0 7183 5 1 1 3258
0 7184 6 1 2 3259 6977
0 7185 5 1 1 3260
0 7186 6 1 2 3261 6978
0 7187 7 1 3 3237 1167 1669
0 7188 7 1 3 3235 1168 1670
0 7189 7 1 3 3233 1169 1671
0 7190 3 5 3 4956 7146 3781
0 7196 7 1 3 3249 1183 1692
0 7197 7 1 3 3247 1184 1693
0 7198 3 5 3 4960 7147 3786
0 7204 6 1 2 3262 7149
0 7205 5 1 1 3263
0 7206 6 1 2 3162 7150
0 7207 7 1 3 3231 1195 1713
0 7208 7 1 3 3245 1208 1736
0 7209 6 2 2 7073 7152
0 7212 6 2 2 7075 7153
0 7215 5 1 1 3252
0 7216 6 1 2 3253 7079
0 7217 5 1 1 3254
0 7218 6 1 2 3255 7083
0 7219 6 2 2 7085 7158
0 7222 6 2 2 7087 7159
0 7225 6 2 2 7089 7160
0 7228 5 1 1 3256
0 7229 6 1 2 3257 7093
0 7236 3 2 2 7173 7125
0 7239 3 2 2 7174 7126
0 7242 3 2 2 7175 7127
0 7245 3 2 2 7176 7040
0 7250 3 6 2 7178 7139
0 7257 3 2 2 7179 7140
0 7260 3 2 2 7180 7141
0 7263 3 2 2 7181 7064
0 7268 6 1 2 3166 7183
0 7269 6 1 2 3168 7185
0 7270 3 5 3 4957 7187 3782
0 7276 3 5 3 4958 7188 3783
0 7282 3 5 3 4959 7189 3784
0 7288 3 5 3 4961 7196 3787
0 7294 3 5 3 3998 7197 3788
0 7300 6 1 2 3223 7205
0 7301 6 2 2 7206 7151
0 7304 3 5 3 4980 7207 3800
0 7310 3 5 3 4984 7208 3805
0 7320 6 1 2 3204 7215
0 7321 6 1 2 3206 7217
0 7328 6 1 2 3214 7228
0 7338 7 1 3 3264 710 1379
0 7339 7 1 3 3269 1372 1380
0 7340 7 1 3 3265 764 1447
0 7341 7 1 3 3270 1442 1448
0 7342 7 1 3 3266 838 1470
0 7349 7 1 3 3271 1464 1471
0 7357 7 1 3 3272 1488 1494
3 7363 5 0 1 3273
0 7364 7 1 3 3267 860 1496
3 7365 5 0 1 3268
0 7394 6 2 2 7268 7184
0 7397 6 2 2 7269 7186
0 7402 6 2 2 7204 7300
0 7405 5 1 1 3274
0 7406 6 1 2 3275 6884
0 7407 5 1 1 3276
0 7408 6 1 2 3277 6888
0 7409 6 2 2 7320 7216
0 7412 6 2 2 7321 7218
0 7415 5 1 1 3278
0 7416 6 1 2 3279 6904
0 7417 5 1 1 3280
0 7418 6 1 2 3281 6908
0 7419 5 1 1 3282
0 7420 6 1 2 3283 6913
0 7421 6 2 2 7328 7229
0 7424 5 1 1 3290
0 7425 5 1 1 3288
0 7426 5 1 1 3286
0 7427 5 1 1 3284
0 7428 5 1 1 3302
0 7429 5 1 1 3300
0 7430 5 1 1 3298
0 7431 5 1 1 3292
3 7432 5 0 1 3293
0 7433 7 1 3 3336 1344 1349
0 7434 7 1 3 3331 687 1350
0 7435 3 1 4 7011 7338 3621 2591
0 7436 7 1 3 3304 711 1382
0 7437 7 1 3 3319 1373 1383
0 7438 7 1 3 3309 712 1385
0 7439 7 1 3 3324 1374 1386
0 7440 7 1 3 3314 713 1388
0 7441 7 1 3 3337 1408 1413
0 7442 7 1 3 3332 742 1414
0 7443 3 1 4 7012 7340 3632 2600
0 7444 7 1 3 3305 765 1449
0 7445 7 1 3 3320 1443 1450
0 7446 7 1 3 3310 766 1451
0 7447 7 1 3 3325 1444 1452
0 7448 7 1 3 3315 767 1453
3 7449 3 0 4 7013 7342 3641 2605
0 7450 7 1 3 3338 1589 1595
0 7451 7 1 3 3333 1090 1596
0 7452 7 1 3 3326 1465 1472
0 7453 7 1 3 3316 839 1473
0 7454 7 1 3 3321 1466 1474
0 7455 7 1 3 3311 840 1476
0 7456 7 1 3 3306 841 1477
0 7457 7 1 3 3339 1626 1634
0 7458 7 1 3 3334 1122 1635
0 7459 7 1 3 3327 1489 1497
0 7460 7 1 3 3317 861 1499
0 7461 7 1 3 3322 1490 1500
0 7462 7 1 3 3312 862 1502
0 7463 7 1 3 3307 863 1503
0 7464 7 1 3 3294 606 602
3 7465 5 0 1 3340
3 7466 5 0 1 3328
3 7467 5 0 1 3323
0 7468 5 1 1 3329
3 7469 3 0 4 7016 7364 3660 2626
3 7470 5 0 1 3335
3 7471 5 0 1 3318
3 7472 5 0 1 3313
3 7473 5 0 1 3308
3 7474 9 0 1 3341
3 7476 9 0 1 3343
0 7479 7 1 2 3330 1616
0 7481 7 1 3 3291 1196 1714
0 7482 7 1 3 3289 1198 1715
0 7483 7 1 3 3287 1199 1716
0 7484 7 1 3 3285 1200 1717
0 7485 7 1 3 3303 1210 1737
0 7486 7 1 3 3301 1211 1738
0 7487 7 1 3 3299 1212 1739
0 7488 7 1 3 3295 1214 1740
0 7489 6 2 2 3220 3296
0 7492 6 1 2 3112 7405
0 7493 6 1 2 3114 7407
0 7498 6 1 2 3140 7415
0 7499 6 1 2 3149 7417
0 7500 6 1 2 3153 7419
3 7503 7 0 9 7105 7166 7167 7168 7169 7424 7425 7426 7427
3 7504 7 0 9 6640 7110 7170 7171 7172 7428 7429 7430 7431
0 7505 3 1 4 7433 7434 3616 2585
3 7506 7 0 2 7435 1360
0 7507 3 1 4 7339 7436 3622 2592
0 7508 3 1 4 7437 7438 3623 2593
0 7509 3 1 4 7439 7440 3624 2594
0 7510 3 1 4 7441 7442 3627 2595
3 7511 7 0 2 7443 1428
0 7512 3 1 4 7341 7444 3633 2601
0 7513 3 1 4 7445 7446 3634 2602
0 7514 3 1 4 7447 7448 3635 2603
3 7515 3 0 4 7450 7451 3646 2610
3 7516 3 0 4 7452 7453 3647 2611
3 7517 3 0 4 7454 7455 3648 2612
3 7518 3 0 4 7349 7456 3649 2613
3 7519 3 0 4 7457 7458 3654 2618
3 7520 3 0 4 7459 7460 3655 2619
3 7521 3 0 4 7461 7462 3656 2620
3 7522 3 0 4 7357 7463 3657 2621
0 7525 3 1 4 4741 7114 2624 7464
0 7526 7 1 3 7468 1684 1694
0 7527 5 1 1 3342
0 7528 5 1 1 3344
0 7529 5 1 1 3345
0 7530 7 1 2 3346 1617
0 7531 3 5 3 4981 7481 3801
0 7537 3 5 3 4982 7482 3802
0 7543 3 5 3 4983 7483 3803
0 7549 3 5 3 5165 7484 3804
0 7555 3 5 3 4985 7485 3806
0 7561 3 5 3 4986 7486 3807
0 7567 3 5 3 4547 7487 3808
0 7573 3 5 3 4987 7488 3809
0 7579 6 2 2 7492 7406
0 7582 6 2 2 7493 7408
0 7585 5 1 1 3347
0 7586 6 1 2 3348 6894
0 7587 5 1 1 3349
0 7588 6 1 2 3350 6900
0 7589 6 2 2 7498 7416
0 7592 6 2 2 7499 7418
0 7595 6 2 2 7500 7420
0 7598 5 1 1 3351
0 7599 6 1 2 3352 6919
3 7600 7 0 2 7505 1333
3 7601 7 0 2 7507 1361
3 7602 7 0 2 7508 1362
3 7603 7 0 2 7509 1364
3 7604 7 0 2 7510 1398
3 7605 7 0 2 7512 1429
3 7606 7 0 2 7513 1431
3 7607 7 0 2 7514 1432
0 7624 7 1 2 3221 3353
0 7625 7 1 2 3354 3297
3 7626 7 0 2 1149 7525
0 7631 7 1 5 565 7527 7528 6805 6930
0 7636 7 1 3 7529 1662 1672
0 7657 6 1 2 3118 7585
0 7658 6 1 2 3123 7587
0 7665 6 1 2 3157 7598
0 7666 7 1 3 3379 1345 1352
0 7667 7 1 3 3355 688 1353
0 7668 7 1 3 3384 1346 1354
0 7669 7 1 3 3364 689 1355
0 7670 7 1 3 3389 1347 1356
0 7671 7 1 3 3369 690 1357
0 7672 7 1 3 3394 1348 1358
0 7673 7 1 3 3374 691 1359
0 7674 7 1 3 3380 1409 1416
0 7675 7 1 3 3356 743 1417
0 7676 7 1 3 3385 1410 1419
0 7677 7 1 3 3365 744 1420
0 7678 7 1 3 3390 1411 1422
0 7679 7 1 3 3370 745 1423
0 7680 7 1 3 3395 1412 1425
0 7681 7 1 3 3375 746 1426
0 7682 7 1 3 3396 1628 1637
0 7683 7 1 3 3376 1123 1638
0 7684 7 1 3 3397 1590 1598
0 7685 7 1 3 3377 1091 1599
0 7686 7 1 3 3391 1591 1601
0 7687 7 1 3 3371 1093 1602
0 7688 7 1 3 3386 1592 1604
0 7689 7 1 3 3366 1094 1605
0 7690 7 1 3 3381 1593 1607
0 7691 7 1 3 3361 1095 1608
0 7692 7 1 3 3392 1629 1640
0 7693 7 1 3 3372 1124 1641
0 7694 7 1 3 3387 1631 1643
0 7695 7 1 3 3367 1125 1644
0 7696 7 1 3 3382 1632 1646
0 7697 7 1 3 3362 1126 1647
3 7698 3 0 2 7624 7625
3 7699 5 0 1 3398
3 7700 5 0 1 3393
3 7701 5 0 1 3388
3 7702 5 0 1 3383
3 7703 7 0 3 1156 7631 247
3 7704 5 0 1 3378
3 7705 5 0 1 3373
3 7706 5 0 1 3368
3 7707 5 0 1 3363
0 7708 5 1 1 3399
0 7709 6 1 2 3400 6739
0 7710 5 1 1 3417
0 7711 6 1 2 3418 6744
0 7712 6 2 2 7657 7586
0 7715 6 2 2 7658 7588
0 7718 5 1 1 3419
0 7719 6 1 2 3420 6772
0 7720 5 1 1 3421
0 7721 6 1 2 3422 6776
0 7722 5 1 1 3423
0 7723 6 1 2 3424 5733
0 7724 6 2 2 7665 7599
0 7727 3 1 4 7666 7667 3617 2586
0 7728 3 1 4 7668 7669 3618 2587
0 7729 3 1 4 7670 7671 3619 2588
0 7730 3 1 4 7672 7673 3620 2589
0 7731 3 1 4 7674 7675 3628 2596
0 7732 3 1 4 7676 7677 3629 2597
0 7733 3 1 4 7678 7679 3630 2598
0 7734 3 1 4 7680 7681 3631 2599
3 7735 3 0 4 7682 7683 3638 2604
3 7736 3 0 4 7684 7685 3642 2606
3 7737 3 0 4 7686 7687 3643 2607
3 7738 3 0 4 7688 7689 3644 2608
3 7739 3 0 4 7690 7691 3645 2609
3 7740 3 0 4 7692 7693 3651 2615
3 7741 3 0 4 7694 7695 3652 2616
3 7742 3 0 4 7696 7697 3653 2617
0 7743 6 1 2 2880 7708
0 7744 6 1 2 2889 7710
0 7749 6 1 2 3043 7718
0 7750 6 1 2 3047 7720
0 7751 6 1 2 2340 7722
3 7754 7 0 2 7727 1334
3 7755 7 0 2 7728 1335
3 7756 7 0 2 7729 1336
3 7757 7 0 2 7730 1337
3 7758 7 0 2 7731 1399
3 7759 7 0 2 7732 1400
3 7760 7 0 2 7733 1401
3 7761 7 0 2 7734 1402
0 7762 6 2 2 7743 7709
0 7765 6 2 2 7744 7711
0 7768 5 1 1 3425
0 7769 6 1 2 3426 6751
0 7770 5 1 1 3427
0 7771 6 1 2 3428 6760
0 7772 6 2 2 7749 7719
0 7775 6 2 2 7750 7721
0 7778 6 2 2 7751 7723
0 7781 5 1 1 3429
0 7782 6 1 2 3430 5735
0 7787 6 1 2 2898 7768
0 7788 6 1 2 2953 7770
0 7795 6 1 2 2344 7781
0 7796 5 1 1 3431
0 7797 6 1 2 3432 6740
0 7798 5 1 1 3433
0 7799 6 1 2 3434 6745
0 7800 6 2 2 7787 7769
0 7803 6 2 2 7788 7771
0 7806 5 1 1 3435
0 7807 6 1 2 3436 6773
0 7808 5 1 1 3437
0 7809 6 1 2 3438 6777
0 7810 5 1 1 3439
0 7811 6 1 2 3440 6782
0 7812 6 2 2 7795 7782
0 7815 6 1 2 2883 7796
0 7816 6 1 2 2892 7798
0 7821 6 1 2 3045 7806
0 7822 6 1 2 3049 7808
0 7823 6 1 2 3051 7810
0 7826 6 2 2 7815 7797
0 7829 6 2 2 7816 7799
0 7832 5 1 1 3441
0 7833 6 1 2 3442 6752
0 7834 5 1 1 3443
0 7835 6 1 2 3457 6761
0 7836 6 2 2 7821 7807
0 7839 6 2 2 7822 7809
0 7842 6 2 2 7823 7811
0 7845 5 1 1 3458
0 7846 6 1 2 3467 6790
0 7851 6 1 2 2900 7832
0 7852 6 1 2 2966 7834
0 7859 6 1 2 3058 7845
0 7860 5 1 1 3468
0 7861 6 1 2 3469 6741
0 7862 5 1 1 3470
0 7863 6 1 2 3471 6746
0 7864 6 2 2 7851 7833
0 7867 6 2 2 7852 7835
0 7870 5 1 1 3472
0 7871 6 1 2 3473 5730
0 7872 5 1 1 3474
0 7873 6 1 2 3475 5732
0 7874 5 1 1 3476
0 7875 6 1 2 3477 6783
0 7876 6 2 2 7859 7846
0 7879 6 1 2 2885 7860
0 7880 6 1 2 2894 7862
0 7885 6 1 2 2330 7870
0 7886 6 1 2 2336 7872
0 7887 6 1 2 3054 7874
0 7890 6 2 2 7879 7861
0 7893 6 2 2 7880 7863
0 7896 5 1 1 3478
0 7897 6 1 2 3479 6753
0 7898 5 1 1 3480
0 7899 6 1 2 3494 6762
0 7900 6 2 2 7885 7871
0 7903 6 2 2 7886 7873
0 7906 6 2 2 7887 7875
0 7909 5 1 1 3495
0 7910 6 1 2 3496 6791
0 7917 6 1 2 2944 7896
0 7918 6 1 2 2968 7898
0 7923 6 1 2 3060 7909
0 7924 5 1 1 3497
0 7925 6 1 2 3498 6680
0 7926 5 1 1 3499
0 7927 6 1 2 3500 6681
0 7928 5 1 1 3501
0 7929 6 1 2 3516 5690
0 7930 5 1 1 3517
0 7931 6 1 2 3518 5691
0 7932 6 2 2 7917 7897
0 7935 6 2 2 7918 7899
0 7938 5 1 1 3519
0 7939 6 1 2 3520 6784
0 7940 6 2 2 7923 7910
0 7943 6 1 2 2887 7924
0 7944 6 1 2 2896 7926
0 7945 6 1 2 2332 7928
0 7946 6 1 2 2338 7930
0 7951 6 1 2 3056 7938
0 7954 6 2 2 7943 7925
0 7957 6 2 2 7944 7927
0 7960 6 2 2 7945 7929
0 7963 6 2 2 7946 7931
0 7966 5 1 1 3521
0 7967 6 1 2 3522 6754
0 7968 5 1 1 3523
0 7969 6 1 2 3524 6755
0 7970 6 2 2 7951 7939
0 7973 5 1 1 3525
0 7974 6 1 2 3526 6785
0 7984 6 1 2 2946 7966
0 7985 6 1 2 3002 7968
0 7987 6 1 2 3062 7973
0 7988 7 1 3 3529 3176 678
0 7989 7 1 3 3527 3076 679
0 7990 7 1 3 3530 3239 568
0 7991 7 1 3 3528 7177 569
0 7992 5 1 1 3535
0 7993 6 1 2 3536 6448
0 7994 7 1 3 3533 3184 733
0 7995 7 1 3 3531 3085 734
0 7996 7 1 3 3534 3251 585
0 7997 7 1 3 3532 7182 586
0 7998 6 2 2 7984 7967
0 8001 6 2 2 7985 7969
0 8004 6 2 2 7987 7974
0 8009 6 1 2 2770 7992
0 8013 3 2 4 7988 7989 7990 7991
0 8017 3 2 4 7994 7995 7996 7997
0 8020 5 1 1 3537
0 8021 6 1 2 3538 6682
0 8022 5 1 1 3539
0 8023 6 1 2 3540 6683
0 8025 6 1 2 8009 7993
0 8026 5 1 1 3541
0 8027 6 1 2 3542 6449
0 8031 6 1 2 2949 8020
0 8032 6 1 2 2951 8022
0 8033 5 1 1 3543
0 8034 6 1 2 2772 8026
0 8035 7 1 2 587 8025
0 8036 5 1 1 3545
0 8037 6 1 2 8031 8021
0 8038 6 1 2 8032 8023
0 8039 6 1 2 8034 8027
0 8040 5 1 1 8038
0 8041 7 1 2 570 8037
0 8042 5 1 1 8039
0 8043 7 1 2 8040 680
0 8044 7 1 2 8042 735
0 8045 3 2 2 8043 8041
0 8048 3 2 2 8044 8035
0 8055 6 1 2 3547 8033
0 8056 5 1 1 3548
0 8057 6 1 2 3549 8036
0 8058 5 1 1 3550
0 8059 6 1 2 3544 8056
0 8060 6 1 2 3546 8058
0 8061 6 2 2 8055 8059
0 8064 6 2 2 8057 8060
0 8071 7 1 3 3553 1186 1695
0 8072 7 1 3 3551 1170 1673
0 8073 5 1 1 3552
0 8074 5 1 1 3554
3 8075 3 0 4 7526 8071 3659 2625
3 8076 3 0 4 7636 8072 3661 2627
0 8077 7 1 2 8073 1114
0 8078 7 1 2 8074 1115
0 8079 3 2 2 7530 8077
0 8082 3 2 2 7479 8078
0 8089 7 1 2 3555 1610
0 8090 7 1 2 3557 1611
0 8091 7 1 2 3556 1613
0 8092 7 1 2 3564 1614
0 8093 3 2 2 8089 3071
0 8096 3 2 2 8090 3072
0 8099 3 2 2 8091 3073
0 8102 3 2 2 8092 3074
0 8113 7 1 3 3571 1467 1478
0 8114 7 1 3 3569 842 1480
0 8115 7 1 3 3572 1491 1505
0 8116 7 1 3 3570 864 1506
0 8117 7 1 3 3567 1376 1389
0 8118 7 1 3 3565 714 1391
0 8119 7 1 3 3568 1445 1454
0 8120 7 1 3 3566 768 1456
0 8121 3 1 4 8117 8118 3662 2703
0 8122 3 1 4 8119 8120 3663 2778
3 8123 3 0 4 8113 8114 3650 2614
3 8124 3 0 4 8115 8116 3658 2622
0 8125 7 1 2 8121 1365
0 8126 7 1 2 8122 1434
3 8127 5 0 1 8125
3 8128 5 0 1 8126
2 2 1 1
2 3 1 1
2 5 1 4
2 6 1 4
2 7 1 4
2 8 1 4
2 9 1 4
2 10 1 4
2 12 1 11
2 13 1 11
2 15 1 14
2 16 1 14
2 18 1 17
2 19 1 17
2 21 1 20
2 22 1 20
2 28 1 27
2 29 1 27
2 30 1 27
2 32 1 31
2 33 1 31
2 35 1 34
2 36 1 34
2 38 1 37
2 39 1 37
2 41 1 40
2 42 1 40
2 44 1 43
2 45 1 43
2 47 1 46
2 48 1 46
2 50 1 49
2 51 1 49
2 55 1 54
2 56 1 54
2 57 1 54
2 58 1 54
2 59 1 54
2 60 1 54
2 62 1 61
2 63 1 61
2 65 1 64
2 66 1 64
2 68 1 67
2 69 1 67
2 71 1 70
2 72 1 70
2 74 1 73
2 75 1 73
2 77 1 76
2 78 1 76
2 84 1 83
2 85 1 83
2 89 1 88
2 90 1 88
2 92 1 91
2 93 1 91
2 95 1 94
2 96 1 94
2 98 1 97
2 99 1 97
2 101 1 100
2 102 1 100
2 104 1 103
2 105 1 103
2 107 1 106
2 108 1 106
2 110 1 109
2 111 1 109
2 124 1 123
2 125 1 123
2 133 1 132
2 134 1 132
2 138 1 137
2 139 1 137
2 142 1 141
2 143 1 141
2 144 1 141
2 147 1 146
2 148 1 146
2 150 1 149
2 151 1 149
2 153 1 152
2 154 1 152
2 156 1 155
2 157 1 155
2 159 1 158
2 160 1 158
2 162 1 161
2 163 1 161
2 165 1 164
2 166 1 164
2 168 1 167
2 169 1 167
2 171 1 170
2 172 1 170
2 174 1 173
2 175 1 173
2 177 1 176
2 178 1 176
2 180 1 179
2 181 1 179
2 183 1 182
2 184 1 182
2 186 1 185
2 187 1 185
2 189 1 188
2 190 1 188
2 192 1 191
2 193 1 191
2 195 1 194
2 196 1 194
2 198 1 197
2 199 1 197
2 201 1 200
2 202 1 200
2 204 1 203
2 205 1 203
2 207 1 206
2 208 1 206
2 211 1 210
2 212 1 210
2 213 1 210
2 214 1 210
2 215 1 210
2 216 1 210
2 219 1 218
2 220 1 218
2 221 1 218
2 222 1 218
2 223 1 218
2 224 1 218
2 227 1 226
2 228 1 226
2 229 1 226
2 230 1 226
2 231 1 226
2 232 1 226
2 235 1 234
2 236 1 234
2 237 1 234
2 238 1 234
2 239 1 234
2 240 1 234
2 243 1 242
2 244 1 242
2 246 1 245
2 247 1 245
2 249 1 248
2 250 1 248
2 252 1 251
2 253 1 251
2 255 1 254
2 256 1 254
2 258 1 257
2 259 1 257
2 260 1 257
2 261 1 257
2 262 1 257
2 263 1 257
2 266 1 265
2 267 1 265
2 268 1 265
2 269 1 265
2 270 1 265
2 271 1 265
2 274 1 273
2 275 1 273
2 276 1 273
2 277 1 273
2 278 1 273
2 279 1 273
2 282 1 281
2 283 1 281
2 284 1 281
2 285 1 281
2 286 1 281
2 287 1 281
2 290 1 289
2 291 1 289
2 294 1 293
2 295 1 293
2 296 1 293
2 297 1 293
2 298 1 293
2 300 1 299
2 301 1 299
2 303 1 302
2 304 1 302
2 305 1 302
2 306 1 302
2 309 1 308
2 310 1 308
2 311 1 308
2 312 1 308
2 313 1 308
2 314 1 308
2 317 1 316
2 318 1 316
2 319 1 316
2 320 1 316
2 321 1 316
2 322 1 316
2 325 1 324
2 326 1 324
2 327 1 324
2 328 1 324
2 329 1 324
2 330 1 324
2 333 1 332
2 334 1 332
2 336 1 335
2 337 1 335
2 339 1 338
2 340 1 338
2 342 1 341
2 343 1 341
2 344 1 341
2 345 1 341
2 346 1 341
2 347 1 341
2 349 1 348
2 350 1 348
2 352 1 351
2 353 1 351
2 354 1 351
2 355 1 351
2 356 1 351
2 357 1 351
2 359 1 358
2 360 1 358
2 362 1 361
2 363 1 361
2 364 1 361
2 365 1 361
2 367 1 366
2 368 1 366
2 370 1 369
2 371 1 369
2 375 1 374
2 376 1 374
2 377 1 374
2 378 1 374
2 379 1 374
2 380 1 374
2 381 1 374
2 382 1 374
2 383 1 374
2 384 1 374
2 385 1 374
2 387 1 386
2 388 1 386
2 390 1 389
2 391 1 389
2 392 1 389
2 393 1 389
2 394 1 389
2 395 1 389
2 396 1 389
2 397 1 389
2 398 1 389
2 399 1 389
2 401 1 400
2 402 1 400
2 403 1 400
2 404 1 400
2 405 1 400
2 406 1 400
2 407 1 400
2 408 1 400
2 409 1 400
2 410 1 400
2 412 1 411
2 413 1 411
2 414 1 411
2 415 1 411
2 416 1 411
2 417 1 411
2 418 1 411
2 419 1 411
2 420 1 411
2 421 1 411
2 423 1 422
2 424 1 422
2 425 1 422
2 426 1 422
2 427 1 422
2 428 1 422
2 429 1 422
2 430 1 422
2 431 1 422
2 432 1 422
2 433 1 422
2 434 1 422
2 436 1 435
2 437 1 435
2 438 1 435
2 439 1 435
2 440 1 435
2 441 1 435
2 442 1 435
2 443 1 435
2 444 1 435
2 445 1 435
2 447 1 446
2 448 1 446
2 449 1 446
2 450 1 446
2 451 1 446
2 452 1 446
2 453 1 446
2 454 1 446
2 455 1 446
2 456 1 446
2 458 1 457
2 459 1 457
2 460 1 457
2 461 1 457
2 462 1 457
2 463 1 457
2 464 1 457
2 465 1 457
2 466 1 457
2 467 1 457
2 469 1 468
2 470 1 468
2 471 1 468
2 472 1 468
2 473 1 468
2 474 1 468
2 475 1 468
2 476 1 468
2 477 1 468
2 478 1 468
2 480 1 479
2 481 1 479
2 482 1 479
2 483 1 479
2 484 1 479
2 485 1 479
2 486 1 479
2 487 1 479
2 488 1 479
2 489 1 479
2 491 1 490
2 492 1 490
2 493 1 490
2 494 1 490
2 495 1 490
2 496 1 490
2 497 1 490
2 498 1 490
2 499 1 490
2 500 1 490
2 501 1 490
2 502 1 490
2 504 1 503
2 505 1 503
2 506 1 503
2 507 1 503
2 508 1 503
2 509 1 503
2 510 1 503
2 511 1 503
2 512 1 503
2 513 1 503
2 515 1 514
2 516 1 514
2 517 1 514
2 518 1 514
2 519 1 514
2 520 1 514
2 521 1 514
2 522 1 514
2 524 1 523
2 525 1 523
2 526 1 523
2 527 1 523
2 528 1 523
2 529 1 523
2 530 1 523
2 531 1 523
2 532 1 523
2 533 1 523
2 535 1 534
2 536 1 534
2 537 1 534
2 538 1 534
2 539 1 534
2 540 1 534
2 541 1 534
2 542 1 534
2 543 1 534
2 544 1 534
2 546 1 545
2 547 1 545
2 548 1 545
2 550 1 549
2 551 1 549
2 553 1 552
2 554 1 552
2 555 1 552
2 557 1 556
2 558 1 556
2 560 1 559
2 561 1 559
2 563 1 562
2 564 1 562
2 565 1 562
2 567 1 566
2 568 1 566
2 569 1 566
2 570 1 566
2 572 1 571
2 573 1 571
2 575 1 574
2 576 1 574
2 578 1 577
2 579 1 577
2 581 1 580
2 582 1 580
2 584 1 583
2 585 1 583
2 586 1 583
2 587 1 583
2 589 1 588
2 590 1 588
2 593 1 592
2 594 1 592
2 600 1 599
2 601 1 599
2 602 1 599
2 604 1 603
2 605 1 603
2 606 1 603
2 608 1 607
2 609 1 607
2 611 1 610
2 612 1 610
2 614 1 613
2 615 1 613
2 617 1 616
2 618 1 616
2 620 1 619
2 621 1 619
2 622 1 619
2 623 1 619
2 624 1 619
2 626 1 625
2 627 1 625
2 628 1 625
2 629 1 625
2 630 1 625
2 632 1 1067
2 633 1 1067
2 634 1 1067
2 635 1 1067
2 636 1 1067
2 637 1 1067
2 638 1 1067
2 639 1 1067
2 640 1 1067
2 641 1 1067
2 642 1 1067
2 643 1 1067
2 644 1 1080
2 645 1 1080
2 646 1 1080
2 647 1 1080
2 648 1 1080
2 649 1 1080
2 650 1 1080
2 651 1 1080
2 652 1 1080
2 653 1 1080
2 654 1 1080
2 655 1 1092
2 656 1 1092
2 657 1 1092
2 658 1 1092
2 659 1 1092
2 660 1 1092
2 661 1 1092
2 662 1 1092
2 663 1 1092
2 664 1 1092
2 665 1 1092
2 666 1 1104
2 667 1 1104
2 668 1 1104
2 669 1 1104
2 670 1 1104
2 671 1 1104
2 672 1 1104
2 673 1 1104
2 674 1 1104
2 675 1 1104
2 676 1 1104
2 677 1 1104
2 678 1 1157
2 679 1 1157
2 680 1 1157
2 681 1 1161
2 682 1 1161
2 683 1 1161
2 684 1 1161
2 685 1 1161
2 686 1 1161
2 687 1 1161
2 688 1 1161
2 689 1 1161
2 690 1 1161
2 691 1 1161
2 692 1 1173
2 693 1 1173
2 694 1 1173
2 695 1 1173
2 696 1 1173
2 697 1 1173
2 698 1 1173
2 699 1 1173
2 700 1 1173
2 701 1 1173
2 702 1 1173
2 703 1 1185
2 704 1 1185
2 705 1 1185
2 706 1 1185
2 707 1 1185
2 708 1 1185
2 710 1 1185
2 711 1 1185
2 712 1 1185
2 713 1 1185
2 714 1 1185
2 715 1 1197
2 716 1 1197
2 717 1 1197
2 718 1 1197
2 719 1 1197
2 720 1 1197
2 721 1 1197
2 722 1 1197
2 723 1 1197
2 724 1 1197
2 725 1 1197
2 726 1 1209
2 727 1 1209
2 728 1 1209
2 729 1 1213
2 730 1 1213
2 731 1 1216
2 732 1 1216
2 733 1 1219
2 734 1 1219
2 735 1 1219
2 736 1 1223
2 737 1 1223
2 738 1 1223
2 739 1 1223
2 740 1 1223
2 741 1 1223
2 742 1 1223
2 743 1 1223
2 744 1 1223
2 745 1 1223
2 746 1 1223
2 747 1 1235
2 748 1 1235
2 749 1 1235
2 750 1 1235
2 751 1 1235
2 752 1 1235
2 753 1 1235
2 754 1 1235
2 755 1 1235
2 756 1 1235
2 757 1 1235
2 758 1 1247
2 759 1 1247
2 760 1 1247
2 761 1 1247
2 762 1 1247
2 763 1 1247
2 764 1 1247
2 765 1 1247
2 766 1 1247
2 767 1 1247
2 768 1 1247
2 769 1 1259
2 770 1 1259
2 771 1 1259
2 772 1 1259
2 773 1 1259
2 774 1 1259
2 775 1 1259
2 776 1 1259
2 777 1 1259
2 778 1 1259
2 779 1 1259
2 780 1 1271
2 781 1 1271
2 782 1 1271
2 783 1 1271
2 784 1 1271
2 785 1 1271
2 786 1 1271
2 787 1 1271
2 788 1 1280
2 789 1 1280
2 790 1 1280
2 791 1 1280
2 792 1 1280
2 793 1 1280
2 794 1 1280
2 795 1 1280
2 796 1 1280
2 797 1 1280
2 798 1 1280
2 799 1 1292
2 800 1 1292
2 801 1 1292
2 802 1 1292
2 803 1 1292
2 804 1 1292
2 805 1 1292
2 806 1 1292
2 807 1 1292
2 808 1 1292
2 809 1 1303
2 810 1 1303
2 811 1 1303
2 812 1 1303
2 813 1 1303
2 814 1 1303
2 815 1 1303
2 817 1 1303
2 818 1 1303
2 819 1 1303
2 820 1 1303
2 821 1 1315
2 822 1 1315
2 823 1 1315
2 824 1 1315
2 825 1 1315
2 826 1 1315
2 827 1 1315
2 828 1 1315
2 829 1 1315
2 830 1 1315
2 831 1 1315
2 832 1 1327
2 833 1 1327
2 834 1 1327
2 835 1 1327
2 836 1 1327
2 837 1 1327
2 838 1 1327
2 839 1 1327
2 840 1 1327
2 841 1 1327
2 842 1 1327
2 843 1 1339
2 844 1 1339
2 845 1 1339
2 846 1 1339
2 847 1 1339
2 848 1 1339
2 849 1 1339
2 850 1 1339
2 851 1 1339
2 852 1 1339
2 853 1 1339
2 854 1 1351
2 855 1 1351
2 856 1 1351
2 857 1 1351
2 858 1 1351
2 859 1 1351
2 860 1 1351
2 861 1 1351
2 862 1 1351
2 863 1 1351
2 864 1 1351
2 865 1 1363
2 866 1 1363
2 867 1 1363
2 868 1 1363
2 869 1 1363
2 870 1 1363
2 871 1 1363
2 872 1 1363
2 873 1 1363
2 874 1 1363
2 875 1 1363
2 876 1 1375
2 877 1 1375
2 878 1 1378
2 879 1 1378
2 880 1 1381
2 881 1 1381
2 882 1 1384
2 883 1 1384
2 884 1 1387
2 885 1 1387
2 886 1 1390
2 887 1 1390
2 888 1 1393
2 889 1 1393
2 890 1 1396
2 891 1 1396
2 892 1 1415
2 893 1 1415
2 894 1 1418
2 895 1 1418
2 896 1 1421
2 897 1 1421
2 898 1 1424
2 899 1 1424
2 900 1 1427
2 901 1 1427
2 902 1 1430
2 903 1 1430
2 904 1 1433
2 905 1 1433
2 906 1 1436
2 907 1 1436
2 908 1 1455
2 909 1 1455
2 910 1 1455
2 911 1 1455
2 912 1 1455
2 913 1 1455
2 914 1 1462
2 915 1 1462
2 916 1 1462
2 917 1 1462
2 918 1 1462
2 919 1 1462
2 920 1 1469
2 921 1 1469
2 922 1 1469
2 923 1 1469
2 924 1 1469
2 925 1 1475
2 926 1 1475
2 927 1 1475
2 928 1 1479
2 929 1 1479
2 930 1 1482
2 931 1 1482
2 932 1 1482
2 933 1 1482
2 934 1 1482
2 935 1 1482
2 936 1 1482
2 937 1 1482
2 938 1 1482
2 939 1 1492
2 940 1 1492
2 941 1 1495
2 942 1 1495
2 943 1 1498
2 944 1 1498
2 945 1 1501
2 946 1 1501
2 947 1 1504
2 948 1 1504
2 949 1 1507
2 950 1 1507
2 951 1 1510
2 952 1 1510
2 953 1 1513
2 954 1 1513
2 955 1 1516
2 956 1 1516
2 957 1 1519
2 958 1 1519
2 959 1 1522
2 960 1 1522
2 961 1 1525
2 962 1 1525
2 963 1 1542
2 964 1 1542
2 965 1 1545
2 966 1 1545
2 967 1 1548
2 968 1 1548
2 969 1 1551
2 970 1 1551
2 971 1 1554
2 972 1 1554
2 973 1 1557
2 974 1 1557
2 975 1 1560
2 976 1 1560
2 977 1 1563
2 978 1 1563
2 979 1 1566
2 980 1 1566
2 981 1 1566
2 982 1 1566
2 983 1 1566
2 984 1 1566
2 985 1 1573
2 986 1 1573
2 987 1 1573
2 988 1 1573
2 989 1 1573
2 990 1 1573
2 991 1 1580
2 992 1 1580
2 993 1 1583
2 994 1 1583
2 995 1 1583
2 996 1 1583
2 997 1 1588
2 998 1 1588
2 999 1 1588
2 1000 1 1588
2 1001 1 1588
2 1002 1 1594
2 1003 1 1594
2 1004 1 1597
2 1005 1 1597
2 1006 1 1600
2 1007 1 1600
2 1008 1 1603
2 1009 1 1603
2 1010 1 1606
2 1011 1 1606
2 1012 1 1609
2 1013 1 1609
2 1014 1 1612
2 1015 1 1612
2 1016 1 1615
2 1017 1 1615
2 1018 1 1618
2 1019 1 1618
2 1020 1 1621
2 1021 1 1621
2 1022 1 1624
2 1023 1 1624
2 1024 1 1627
2 1025 1 1627
2 1026 1 1630
2 1027 1 1630
2 1028 1 1633
2 1029 1 1633
2 1030 1 1636
2 1031 1 1636
2 1032 1 1639
2 1033 1 1639
2 1034 1 1642
2 1035 1 1642
2 1036 1 1645
2 1037 1 1645
2 1038 1 1648
2 1039 1 1648
2 1040 1 1651
2 1041 1 1651
2 1044 1 1654
2 1045 1 1654
2 1046 1 1657
2 1047 1 1657
2 1048 1 1660
2 1049 1 1660
2 1050 1 1663
2 1051 1 1663
2 1052 1 1663
2 1053 1 1663
2 1054 1 1663
2 1055 1 1663
2 1056 1 1663
2 1057 1 1663
2 1058 1 1663
2 1059 1 1663
2 1060 1 1663
2 1061 1 1675
2 1062 1 1675
2 1063 1 1675
2 1064 1 1675
2 1065 1 1675
2 1068 1 1675
2 1069 1 1675
2 1070 1 1675
2 1071 1 1675
2 1072 1 1685
2 1073 1 1685
2 1074 1 1685
2 1075 1 1685
2 1076 1 1685
2 1077 1 1685
2 1078 1 1685
2 1079 1 1685
2 1081 1 1685
2 1082 1 1685
2 1083 1 1685
2 1084 1 1697
2 1085 1 1697
2 1086 1 1697
2 1087 1 1697
2 1088 1 1697
2 1089 1 1697
2 1090 1 1697
2 1091 1 1697
2 1093 1 1697
2 1094 1 1697
2 1095 1 1697
2 1096 1 1709
2 1097 1 1709
2 1098 1 1709
2 1099 1 1709
2 1100 1 1709
2 1101 1 1709
2 1102 1 1709
2 1103 1 1709
2 1105 1 1709
2 1106 1 1709
2 1107 1 1709
2 1108 1 1721
2 1109 1 1721
2 1110 1 1721
2 1111 1 1721
2 1112 1 1721
2 1113 1 1727
2 1114 1 1727
2 1115 1 1727
2 1116 1 1731
2 1117 1 1731
2 1118 1 1731
2 1119 1 1731
2 1120 1 1731
2 1121 1 1731
2 1122 1 1731
2 1123 1 1731
2 1124 1 1731
2 1125 1 1731
2 1126 1 1731
2 1127 1 1743
2 1128 1 1743
2 1129 1 1743
2 1130 1 1743
2 1131 1 1743
2 1132 1 1743
2 1133 1 1743
2 1134 1 1743
2 1135 1 1743
2 1136 1 1743
2 1158 1 1743
2 1159 1 1755
2 1160 1 1755
2 1162 1 1758
2 1163 1 1758
2 1164 1 1761
2 1165 1 1761
2 1166 1 1761
2 1167 1 1761
2 1168 1 1761
2 1169 1 1761
2 1170 1 1761
2 1171 1 1769
2 1172 1 1769
2 1174 1 1769
2 1175 1 1769
2 1176 1 1769
2 1177 1 1769
2 1178 1 1769
2 1179 1 1777
2 1180 1 1777
2 1181 1 1777
2 1182 1 1777
2 1183 1 1777
2 1184 1 1777
2 1186 1 1777
2 1187 1 1785
2 1188 1 1785
2 1189 1 1785
2 1190 1 1785
2 1191 1 1785
2 1192 1 1785
2 1193 1 1785
2 1194 1 1793
2 1195 1 1793
2 1196 1 1793
2 1198 1 1793
2 1199 1 1793
2 1200 1 1793
2 1201 1 1800
2 1202 1 1800
2 1203 1 1800
2 1204 1 1800
2 1205 1 1800
2 1206 1 1800
2 1207 1 1807
2 1208 1 1807
2 1210 1 1807
2 1211 1 1807
2 1212 1 1807
2 1214 1 1807
2 1215 1 1814
2 1217 1 1814
2 1218 1 1814
2 1220 1 1814
2 1221 1 1814
2 1222 1 1814
2 1224 1 1821
2 1225 1 1821
2 1226 1 1824
2 1227 1 1824
2 1228 1 1827
2 1229 1 1827
2 1230 1 1830
2 1231 1 1830
2 1232 1 1833
2 1233 1 1833
2 1234 1 1836
2 1236 1 1836
2 1237 1 1839
2 1238 1 1839
2 1239 1 1842
2 1240 1 1842
2 1241 1 1845
2 1242 1 1845
2 1243 1 1848
2 1244 1 1848
2 1245 1 1851
2 1246 1 1851
2 1248 1 1854
2 1249 1 1854
2 1250 1 1857
2 1251 1 1857
2 1252 1 1860
2 1253 1 1860
2 1254 1 1863
2 1255 1 1863
2 1256 1 1866
2 1257 1 1866
2 1258 1 1869
2 1260 1 1869
2 1261 1 1872
2 1262 1 1872
2 1263 1 1875
2 1264 1 1875
2 1265 1 1878
2 1266 1 1878
2 1267 1 1881
2 1268 1 1881
2 1269 1 1884
2 1270 1 1884
2 1272 1 1887
2 1273 1 1887
2 1274 1 1890
2 1275 1 1890
2 1276 1 1893
2 1277 1 1893
2 1278 1 1896
2 1279 1 1896
2 1281 1 1899
2 1282 1 1899
2 1283 1 1902
2 1284 1 1902
2 1285 1 1905
2 1286 1 1905
2 1287 1 1908
2 1288 1 1908
2 1289 1 1911
2 1290 1 1911
2 1291 1 1914
2 1293 1 1914
2 1294 1 1917
2 1295 1 1917
2 1296 1 1920
2 1297 1 1920
2 1298 1 1923
2 1299 1 1923
2 1300 1 1926
2 1301 1 1926
2 1302 1 1929
2 1304 1 1929
2 1305 1 1932
2 1306 1 1932
2 1307 1 1935
2 1308 1 1935
2 1309 1 1938
2 1310 1 1938
2 1311 1 1941
2 1312 1 1941
2 1313 1 1944
2 1314 1 1944
2 1316 1 1947
2 1317 1 1947
2 1318 1 1950
2 1319 1 1950
2 1320 1 1953
2 1321 1 1953
2 1322 1 1956
2 1323 1 1956
2 1324 1 1959
2 1325 1 1959
2 1326 1 1962
2 1328 1 1962
2 1329 1 1965
2 1330 1 1965
2 1331 1 1968
2 1332 1 1968
2 1333 1 2647
2 1334 1 2647
2 1335 1 2647
2 1336 1 2647
2 1337 1 2647
2 1338 1 2653
2 1340 1 2653
2 1341 1 2653
2 1342 1 2653
2 1343 1 2653
2 1344 1 2653
2 1345 1 2653
2 1346 1 2653
2 1347 1 2653
2 1348 1 2653
2 1349 1 2664
2 1350 1 2664
2 1352 1 2664
2 1353 1 2664
2 1354 1 2664
2 1355 1 2664
2 1356 1 2664
2 1357 1 2664
2 1358 1 2664
2 1359 1 2664
2 1360 1 2675
2 1361 1 2675
2 1362 1 2675
2 1364 1 2675
2 1365 1 2675
2 1366 1 2681
2 1367 1 2681
2 1368 1 2681
2 1369 1 2681
2 1370 1 2681
2 1371 1 2681
2 1372 1 2681
2 1373 1 2681
2 1374 1 2681
2 1376 1 2681
2 1377 1 2692
2 1379 1 2692
2 1380 1 2692
2 1382 1 2692
2 1383 1 2692
2 1385 1 2692
2 1386 1 2692
2 1388 1 2692
2 1389 1 2692
2 1391 1 2692
2 1392 1 2704
2 1394 1 2704
2 1395 1 2704
2 1397 1 2704
2 1398 1 2722
2 1399 1 2722
2 1400 1 2722
2 1401 1 2722
2 1402 1 2722
2 1403 1 2728
2 1404 1 2728
2 1405 1 2728
2 1406 1 2728
2 1407 1 2728
2 1408 1 2728
2 1409 1 2728
2 1410 1 2728
2 1411 1 2728
2 1412 1 2728
2 1413 1 2739
2 1414 1 2739
2 1416 1 2739
2 1417 1 2739
2 1419 1 2739
2 1420 1 2739
2 1422 1 2739
2 1423 1 2739
2 1425 1 2739
2 1426 1 2739
2 1428 1 2750
2 1429 1 2750
2 1431 1 2750
2 1432 1 2750
2 1434 1 2750
2 1435 1 2756
2 1437 1 2756
2 1438 1 2756
2 1439 1 2756
2 1440 1 2756
2 1441 1 2756
2 1442 1 2756
2 1443 1 2756
2 1444 1 2756
2 1445 1 2756
2 1446 1 2767
2 1447 1 2767
2 1448 1 2767
2 1449 1 2767
2 1450 1 2767
2 1451 1 2767
2 1452 1 2767
2 1453 1 2767
2 1454 1 2767
2 1456 1 2767
2 1457 1 2779
2 1458 1 2779
2 1459 1 2779
2 1460 1 2779
2 1461 1 2779
2 1463 1 2779
2 1464 1 2779
2 1465 1 2779
2 1466 1 2779
2 1467 1 2779
2 1468 1 2790
2 1470 1 2790
2 1471 1 2790
2 1472 1 2790
2 1473 1 2790
2 1474 1 2790
2 1476 1 2790
2 1477 1 2790
2 1478 1 2790
2 1480 1 2790
2 1481 1 2801
2 1483 1 2801
2 1484 1 2801
2 1485 1 2801
2 1486 1 2801
2 1487 1 2801
2 1488 1 2801
2 1489 1 2801
2 1490 1 2801
2 1491 1 2801
2 1493 1 2812
2 1494 1 2812
2 1496 1 2812
2 1497 1 2812
2 1499 1 2812
2 1500 1 2812
2 1502 1 2812
2 1503 1 2812
2 1505 1 2812
2 1506 1 2812
2 1508 1 2855
2 1509 1 2855
2 1511 1 2855
2 1512 1 2855
2 1514 1 2855
2 1515 1 2861
2 1517 1 2861
2 1518 1 2861
2 1520 1 2861
2 1521 1 2861
2 1523 1 2877
2 1524 1 2877
2 1526 1 2877
2 1527 1 2877
2 1528 1 2882
2 1529 1 2882
2 1530 1 2882
2 1531 1 2882
2 1532 1 2882
2 1533 1 2882
2 1534 1 2882
2 1535 1 2882
2 1536 1 2891
2 1537 1 2891
2 1538 1 2891
2 1539 1 2891
2 1540 1 2891
2 1541 1 2891
2 1543 1 2891
2 1544 1 2891
2 1546 1 2891
2 1547 1 2942
2 1549 1 2942
2 1550 1 2942
2 1552 1 2942
2 1553 1 2942
2 1555 1 2948
2 1556 1 2948
2 1558 1 2948
2 1559 1 2948
2 1561 1 2948
2 1562 1 2964
2 1564 1 2964
2 1565 1 2964
2 1567 1 2964
2 1568 1 3000
2 1569 1 3000
2 1570 1 3003
2 1571 1 3003
2 1572 1 3007
2 1574 1 3007
2 1575 1 3010
2 1576 1 3010
2 1577 1 3035
2 1578 1 3035
2 1579 1 3038
2 1581 1 3038
2 1582 1 3041
2 1584 1 3041
2 1585 1 3041
2 1586 1 3041
2 1587 1 3041
2 1589 1 3041
2 1590 1 3041
2 1591 1 3041
2 1592 1 3041
2 1593 1 3041
2 1595 1 3052
2 1596 1 3052
2 1598 1 3052
2 1599 1 3052
2 1601 1 3052
2 1602 1 3052
2 1604 1 3052
2 1605 1 3052
2 1607 1 3052
2 1608 1 3052
2 1610 1 3063
2 1611 1 3063
2 1613 1 3063
2 1614 1 3063
2 1616 1 3068
2 1617 1 3068
2 1619 1 3075
2 1620 1 3075
2 1622 1 3075
2 1623 1 3075
2 1625 1 3075
2 1626 1 3075
2 1628 1 3075
2 1629 1 3075
2 1631 1 3075
2 1632 1 3075
2 1634 1 3086
2 1635 1 3086
2 1637 1 3086
2 1638 1 3086
2 1640 1 3086
2 1641 1 3086
2 1643 1 3086
2 1644 1 3086
2 1646 1 3086
2 1647 1 3086
2 1649 1 3097
2 1650 1 3097
2 1652 1 3097
2 1653 1 3097
2 1655 1 3097
2 1656 1 3097
2 1658 1 3097
2 1659 1 3097
2 1661 1 3097
2 1662 1 3097
2 1664 1 3108
2 1665 1 3108
2 1666 1 3108
2 1667 1 3108
2 1668 1 3108
2 1669 1 3108
2 1670 1 3108
2 1671 1 3108
2 1672 1 3108
2 1673 1 3108
2 1674 1 3119
2 1676 1 3119
2 1677 1 3119
2 1678 1 3119
2 1679 1 3119
2 1680 1 3119
2 1681 1 3119
2 1682 1 3119
2 1683 1 3119
2 1684 1 3119
2 1686 1 3130
2 1687 1 3130
2 1688 1 3130
2 1689 1 3130
2 1690 1 3130
2 1691 1 3130
2 1692 1 3130
2 1693 1 3130
2 1694 1 3130
2 1695 1 3130
2 1696 1 3147
2 1698 1 3147
2 1699 1 3147
2 1700 1 3147
2 1701 1 3147
2 1702 1 3147
2 1703 1 3147
2 1704 1 3147
2 1705 1 3147
2 1706 1 3147
2 1707 1 3158
2 1708 1 3158
2 1710 1 3158
2 1711 1 3158
2 1712 1 3158
2 1713 1 3158
2 1714 1 3158
2 1715 1 3158
2 1716 1 3158
2 1717 1 3158
2 1718 1 3169
2 1719 1 3169
2 1720 1 3169
2 1722 1 3169
2 1723 1 3169
2 1724 1 3169
2 1725 1 3169
2 1726 1 3169
2 1728 1 3169
2 1729 1 3169
2 1730 1 3180
2 1732 1 3180
2 1733 1 3180
2 1734 1 3180
2 1735 1 3180
2 1736 1 3180
2 1737 1 3180
2 1738 1 3180
2 1739 1 3180
2 1740 1 3180
2 1741 1 3191
2 1742 1 3191
2 1744 1 3200
2 1745 1 3200
2 1746 1 3456
2 1747 1 3456
2 1748 1 3691
2 1749 1 3691
2 1750 1 3691
2 1751 1 3691
2 1752 1 3691
2 1753 1 3691
2 1754 1 3691
2 1756 1 3691
2 1757 1 3705
2 1759 1 3705
2 1760 1 3732
2 1762 1 3732
2 1763 1 3732
2 1764 1 3732
2 1765 1 3732
2 1766 1 3771
2 1767 1 3771
2 1768 1 3771
2 1770 1 3775
2 1771 1 3775
2 1772 1 3775
2 1773 1 3789
2 1774 1 3789
2 1775 1 3789
2 1776 1 3793
2 1778 1 3793
2 1779 1 3793
2 1780 1 3797
2 1781 1 3797
2 1782 1 3810
2 1783 1 3810
2 1784 1 3813
2 1786 1 3813
2 1787 1 3816
2 1788 1 3816
2 1789 1 3819
2 1790 1 3819
2 1791 1 3824
2 1792 1 3824
2 1794 1 3842
2 1795 1 3842
2 1796 1 3842
2 1797 1 3842
2 1798 1 3842
2 1799 1 3842
2 1801 1 3849
2 1802 1 3849
2 1803 1 3849
2 1804 1 3849
2 1805 1 3849
2 1806 1 3855
2 1808 1 3855
2 1809 1 3855
2 1810 1 3855
2 1811 1 3855
2 1812 1 3861
2 1813 1 3861
2 1815 1 3861
2 1816 1 3861
2 1817 1 3861
2 1818 1 3867
2 1819 1 3867
2 1820 1 3867
2 1822 1 3867
2 1823 1 3867
2 1825 1 3873
2 1826 1 3873
2 1828 1 3873
2 1829 1 3873
2 1831 1 3873
2 1832 1 3873
2 1834 1 3873
2 1835 1 3881
2 1837 1 3881
2 1838 1 3881
2 1840 1 3881
2 1841 1 3881
2 1843 1 3887
2 1844 1 3887
2 1846 1 3887
2 1847 1 3887
2 1849 1 3887
2 1850 1 3893
2 1852 1 3893
2 1853 1 3893
2 1855 1 3893
2 1856 1 3893
2 1858 1 3911
2 1859 1 3911
2 1861 1 3921
2 1862 1 3921
2 1864 1 3921
2 1865 1 3921
2 1867 1 3921
2 1868 1 3927
2 1870 1 3927
2 1871 1 3927
2 1873 1 3927
2 1874 1 3927
2 1876 1 3933
2 1877 1 3933
2 1879 1 3933
2 1880 1 3933
2 1882 1 3933
2 1883 1 3942
2 1885 1 3942
2 1886 1 3942
2 1888 1 3942
2 1889 1 3942
2 1891 1 3948
2 1892 1 3948
2 1894 1 3948
2 1895 1 3948
2 1897 1 3948
2 1898 1 3948
2 1900 1 3948
2 1901 1 3956
2 1903 1 3956
2 1904 1 3956
2 1906 1 3956
2 1907 1 3956
2 1909 1 3962
2 1910 1 3962
2 1912 1 3962
2 1913 1 3962
2 1915 1 3962
2 1916 1 3968
2 1918 1 3968
2 1919 1 3968
2 1921 1 3968
2 1922 1 3968
2 1924 1 3968
2 1925 1 3984
2 1927 1 3984
2 1928 1 4008
2 1930 1 4008
2 1931 1 4011
2 1933 1 4011
2 1934 1 4021
2 1936 1 4021
2 1937 1 4067
2 1939 1 4067
2 1940 1 4080
2 1942 1 4080
2 1943 1 4080
2 1945 1 4088
2 1946 1 4088
2 1948 1 4091
2 1949 1 4091
2 1951 1 4094
2 1952 1 4094
2 1954 1 4097
2 1955 1 4097
2 1957 1 4100
2 1958 1 4100
2 1960 1 4103
2 1961 1 4103
2 1963 1 4106
2 1964 1 4106
2 1966 1 4109
2 1967 1 4109
2 1969 1 4144
2 1970 1 4144
2 1971 1 4147
2 1973 1 4147
2 1974 1 4150
2 1975 1 4150
2 1976 1 4153
2 1977 1 4153
2 1978 1 4156
2 1979 1 4156
2 1980 1 4159
2 1981 1 4159
2 1982 1 4188
2 1983 1 4188
2 1984 1 4191
2 1985 1 4191
2 1986 1 4200
2 1987 1 4200
2 1988 1 4203
2 1989 1 4203
2 1990 1 4206
2 1991 1 4206
2 1992 1 4209
2 1993 1 4209
2 1994 1 4212
2 1995 1 4212
2 1996 1 4215
2 1997 1 4215
2 1998 1 4219
2 1999 1 4219
2 2000 1 4225
2 2001 1 4225
2 2002 1 4228
2 2003 1 4228
2 2004 1 4231
2 2005 1 4231
2 2006 1 4234
2 2007 1 4234
2 2008 1 4237
2 2009 1 4237
2 2010 1 4240
2 2011 1 4240
2 2012 1 4243
2 2013 1 4243
2 2014 1 4246
2 2015 1 4246
2 2016 1 4249
2 2017 1 4249
2 2018 1 4252
2 2019 1 4252
2 2020 1 4255
2 2021 1 4255
2 2022 1 4258
2 2023 1 4258
2 2024 1 4264
2 2025 1 4264
2 2026 1 4280
2 2027 1 4280
2 2028 1 4280
2 2029 1 4284
2 2030 1 4284
2 2031 1 4284
2 2032 1 4284
2 2033 1 4284
2 2034 1 4290
2 2035 1 4290
2 2036 1 4290
2 2037 1 4290
2 2038 1 4290
2 2039 1 4290
2 2040 1 4298
2 2041 1 4298
2 2042 1 4301
2 2043 1 4301
2 2044 1 4301
2 2045 1 4305
2 2046 1 4305
2 2047 1 4305
2 2048 1 4305
2 2049 1 4310
2 2050 1 4310
2 2051 1 4310
2 2052 1 4310
2 2053 1 4310
2 2055 1 4316
2 2056 1 4316
2 2057 1 4316
2 2058 1 4320
2 2059 1 4320
2 2062 1 4320
2 2063 1 4320
2 2064 1 4325
2 2065 1 4325
2 2066 1 4325
2 2067 1 4325
2 2068 1 4325
2 2069 1 4332
2 2070 1 4332
2 2071 1 4332
2 2072 1 4336
2 2073 1 4336
2 2074 1 4336
2 2075 1 4336
2 2076 1 4336
2 2077 1 4342
2 2078 1 4342
2 2079 1 4342
2 2080 1 4342
2 2081 1 4342
2 2082 1 4342
2 2083 1 4349
2 2084 1 4349
2 2085 1 4349
2 2086 1 4349
2 2087 1 4349
2 2088 1 4349
2 2089 1 4349
2 2090 1 4357
2 2091 1 4357
2 2092 1 4357
2 2093 1 4357
2 2094 1 4357
2 2095 1 4357
2 2096 1 4364
2 2097 1 4364
2 2098 1 4364
2 2099 1 4364
2 2100 1 4364
2 2101 1 4364
2 2102 1 4364
2 2103 1 4364
2 2104 1 4364
2 2105 1 4364
2 2106 1 4375
2 2107 1 4375
2 2108 1 4375
2 2109 1 4379
2 2110 1 4379
2 2111 1 4379
2 2112 1 4379
2 2113 1 4379
2 2114 1 4385
2 2115 1 4385
2 2116 1 4385
2 2117 1 4385
2 2118 1 4385
2 2119 1 4385
2 2120 1 4396
2 2121 1 4396
2 2122 1 4396
2 2123 1 4400
2 2124 1 4400
2 2125 1 4400
2 2126 1 4400
2 2127 1 4405
2 2128 1 4405
2 2129 1 4405
2 2130 1 4405
2 2131 1 4405
2 2132 1 4405
2 2133 1 4412
2 2134 1 4412
2 2135 1 4412
2 2136 1 4412
2 2137 1 4412
2 2138 1 4418
2 2140 1 4418
2 2141 1 4418
2 2143 1 4418
2 2144 1 4418
2 2145 1 4418
2 2146 1 4425
2 2147 1 4425
2 2148 1 4425
2 2149 1 4425
2 2150 1 4425
2 2151 1 4425
2 2152 1 4425
2 2153 1 4425
2 2154 1 4425
2 2155 1 4425
2 2156 1 4436
2 2157 1 4436
2 2158 1 4436
2 2159 1 4440
2 2160 1 4440
2 2161 1 4440
2 2162 1 4440
2 2163 1 4445
2 2164 1 4445
2 2165 1 4445
2 2166 1 4445
2 2167 1 4445
2 2168 1 4456
2 2169 1 4456
2 2170 1 4456
2 2171 1 4456
2 2172 1 4456
2 2173 1 4462
2 2174 1 4462
2 2175 1 4462
2 2176 1 4462
2 2177 1 4462
2 2178 1 4462
2 2179 1 4469
2 2180 1 4469
2 2181 1 4469
2 2182 1 4469
2 2183 1 4469
2 2184 1 4469
2 2185 1 4469
2 2186 1 4477
2 2187 1 4477
2 2188 1 4477
2 2189 1 4477
2 2190 1 4477
2 2191 1 4477
2 2192 1 4512
2 2193 1 4512
2 2194 1 4524
2 2195 1 4524
2 2196 1 4524
2 2197 1 4532
2 2198 1 4532
2 2199 1 4532
2 2200 1 4548
2 2201 1 4548
2 2202 1 4551
2 2203 1 4551
2 2204 1 4554
2 2205 1 4554
2 2206 1 4557
2 2207 1 4557
2 2208 1 4560
2 2209 1 4560
2 2210 1 4563
2 2211 1 4563
2 2212 1 4566
2 2213 1 4566
2 2214 1 4569
2 2215 1 4569
2 2216 1 4572
2 2217 1 4572
2 2218 1 4575
2 2219 1 4575
2 2220 1 4578
2 2221 1 4578
2 2222 1 4581
2 2223 1 4581
2 2224 1 4584
2 2225 1 4584
2 2226 1 4587
2 2227 1 4587
2 2228 1 4590
2 2229 1 4590
2 2230 1 4593
2 2231 1 4593
2 2232 1 4596
2 2233 1 4596
2 2234 1 4599
2 2235 1 4599
2 2236 1 4602
2 2237 1 4602
2 2238 1 4605
2 2239 1 4605
2 2240 1 4608
2 2241 1 4608
2 2242 1 4611
2 2243 1 4611
2 2244 1 4614
2 2245 1 4614
2 2246 1 4617
2 2247 1 4617
2 2248 1 4621
2 2249 1 4621
2 2250 1 4624
2 2251 1 4624
2 2252 1 4627
2 2253 1 4627
2 2254 1 4630
2 2255 1 4630
2 2256 1 4633
2 2257 1 4633
2 2258 1 4637
2 2259 1 4637
2 2260 1 4640
2 2261 1 4640
2 2262 1 4643
2 2263 1 4643
2 2264 1 4646
2 2265 1 4646
2 2266 1 4649
2 2267 1 4649
2 2268 1 4652
2 2269 1 4652
2 2270 1 4655
2 2271 1 4655
2 2272 1 4658
2 2273 1 4658
2 2274 1 4662
2 2275 1 4662
2 2276 1 4665
2 2277 1 4665
2 2278 1 4668
2 2279 1 4668
2 2280 1 4671
2 2281 1 4671
2 2282 1 4674
2 2283 1 4674
2 2284 1 4677
2 2285 1 4677
2 2286 1 4680
2 2287 1 4680
2 2288 1 4683
2 2289 1 4683
2 2290 1 4686
2 2291 1 4686
2 2292 1 4689
2 2293 1 4689
2 2294 1 4692
2 2295 1 4692
2 2296 1 4695
2 2297 1 4695
2 2298 1 4698
2 2299 1 4698
2 2300 1 4939
2 2301 1 4939
2 2302 1 5049
2 2303 1 5049
2 2304 1 5150
2 2305 1 5150
2 2306 1 5157
2 2307 1 5157
2 2308 1 5166
2 2310 1 5166
2 2311 1 5169
2 2312 1 5169
2 2313 1 5173
2 2314 1 5173
2 2315 1 5177
2 2316 1 5177
2 2317 1 5180
2 2318 1 5180
2 2319 1 5183
2 2320 1 5183
2 2321 1 5186
2 2322 1 5186
2 2323 1 5189
2 2324 1 5189
2 2325 1 5192
2 2326 1 5192
2 2327 1 5195
2 2328 1 5195
2 2329 1 5199
2 2330 1 5199
2 2331 1 5202
2 2332 1 5202
2 2333 1 5205
2 2334 1 5205
2 2335 1 5208
2 2336 1 5208
2 2337 1 5211
2 2338 1 5211
2 2339 1 5214
2 2340 1 5214
2 2341 1 5217
2 2342 1 5217
2 2343 1 5220
2 2344 1 5220
2 2345 1 5236
2 2346 1 5236
2 2347 1 5264
2 2348 1 5264
2 2351 1 5264
2 2352 1 5264
2 2353 1 5264
2 2354 1 5264
2 2355 1 5264
2 2356 1 5264
2 2357 1 5264
2 2358 1 5284
2 2359 1 5284
2 2360 1 5284
2 2361 1 5284
2 2362 1 5284
2 2363 1 5284
2 2364 1 5284
2 2365 1 5284
2 2366 1 5284
2 2367 1 5284
2 2368 1 5284
2 2369 1 5284
2 2370 1 5284
2 2371 1 5315
2 2372 1 5315
2 2373 1 5315
2 2374 1 5319
2 2375 1 5319
2 2376 1 5324
2 2377 1 5324
2 2378 1 5324
2 2379 1 5328
2 2380 1 5328
2 2381 1 5346
2 2382 1 5346
2 2383 1 5371
2 2384 1 5371
2 2385 1 5374
2 2386 1 5374
2 2388 1 5377
2 2389 1 5377
2 2390 1 5382
2 2391 1 5382
2 2392 1 5385
2 2393 1 5385
2 2394 1 5389
2 2395 1 5389
2 2396 1 5389
2 2397 1 5389
2 2398 1 5389
2 2399 1 5389
2 2400 1 5396
2 2401 1 5396
2 2402 1 5396
2 2403 1 5396
2 2404 1 5396
2 2405 1 5396
2 2406 1 5396
2 2407 1 5396
2 2408 1 5396
2 2409 1 5396
2 2410 1 5407
2 2411 1 5407
2 2412 1 5407
2 2413 1 5407
2 2414 1 5407
2 2415 1 5407
2 2416 1 5407
2 2417 1 5407
2 2418 1 5407
2 2419 1 5407
2 2420 1 5418
2 2421 1 5418
2 2422 1 5418
2 2423 1 5418
2 2424 1 5418
2 2425 1 5424
2 2426 1 5424
2 2427 1 5424
2 2428 1 5424
2 2429 1 5424
2 2430 1 5424
2 2431 1 5431
2 2432 1 5431
2 2433 1 5431
2 2434 1 5431
2 2435 1 5431
2 2436 1 5431
2 2437 1 5431
2 2438 1 5431
2 2439 1 5431
2 2440 1 5441
2 2441 1 5441
2 2442 1 5441
2 2443 1 5441
2 2444 1 5441
2 2445 1 5441
2 2446 1 5441
2 2447 1 5441
2 2448 1 5441
2 2449 1 5441
2 2450 1 5452
2 2451 1 5452
2 2452 1 5452
2 2453 1 5452
2 2454 1 5452
2 2455 1 5452
2 2456 1 5452
2 2457 1 5452
2 2458 1 5452
2 2459 1 5462
2 2460 1 5462
2 2461 1 5462
2 2462 1 5462
2 2463 1 5462
2 2464 1 5462
2 2465 1 5470
2 2466 1 5470
2 2467 1 5470
2 2468 1 5470
2 2469 1 5470
2 2470 1 5470
2 2471 1 5477
2 2472 1 5477
2 2473 1 5477
2 2474 1 5477
2 2475 1 5477
2 2476 1 5477
2 2477 1 5477
2 2478 1 5477
2 2479 1 5477
2 2480 1 5477
2 2481 1 5488
2 2482 1 5488
2 2483 1 5488
2 2484 1 5488
2 2485 1 5488
2 2486 1 5488
2 2487 1 5488
2 2488 1 5488
2 2489 1 5488
2 2490 1 5498
2 2491 1 5498
2 2492 1 5498
2 2493 1 5498
2 2494 1 5498
2 2495 1 5498
2 2496 1 5498
2 2497 1 5506
2 2498 1 5506
2 2499 1 5506
2 2500 1 5506
2 2501 1 5506
2 2502 1 5506
2 2503 1 5506
2 2504 1 5506
2 2505 1 5506
2 2506 1 5506
2 2507 1 5506
2 2508 1 5506
2 2509 1 5506
2 2510 1 5520
2 2511 1 5520
2 2512 1 5520
2 2513 1 5520
2 2514 1 5520
2 2515 1 5520
2 2516 1 5520
2 2517 1 5520
2 2518 1 5520
2 2519 1 5520
2 2520 1 5520
2 2521 1 5520
2 2522 1 5520
2 2523 1 5520
2 2524 1 5520
2 2525 1 5536
2 2526 1 5536
2 2528 1 5536
2 2529 1 5536
2 2530 1 5536
2 2531 1 5536
2 2532 1 5536
2 2533 1 5536
2 2534 1 5536
2 2535 1 5536
2 2536 1 5536
2 2537 1 5536
2 2538 1 5549
2 2539 1 5549
2 2540 1 5549
2 2541 1 5549
2 2542 1 5549
2 2543 1 5555
2 2544 1 5555
2 2545 1 5555
2 2546 1 5555
2 2547 1 5555
2 2548 1 5555
2 2549 1 5562
2 2550 1 5562
2 2551 1 5562
2 2552 1 5562
2 2553 1 5562
2 2554 1 5562
2 2555 1 5562
2 2556 1 5562
2 2557 1 5562
2 2558 1 5562
2 2559 1 5573
2 2560 1 5573
2 2561 1 5573
2 2562 1 5573
2 2563 1 5573
2 2564 1 5579
2 2565 1 5579
2 2566 1 5579
2 2567 1 5579
2 2568 1 5579
2 2569 1 5579
2 2570 1 5595
2 2571 1 5595
2 2572 1 5595
2 2573 1 5595
2 2574 1 5595
2 2575 1 5595
2 2576 1 5595
2 2577 1 5595
2 2578 1 5595
2 2579 1 5595
2 2580 1 5606
2 2581 1 5606
2 2582 1 5606
2 2583 1 5606
2 2648 1 5606
2 2649 1 5606
2 2650 1 5606
2 2651 1 5606
2 2652 1 5606
2 2654 1 5624
2 2655 1 5624
2 2656 1 5624
2 2657 1 5624
2 2658 1 5624
2 2659 1 5624
2 2660 1 5624
2 2661 1 5624
2 2662 1 5624
2 2663 1 5634
2 2665 1 5634
2 2666 1 5634
2 2667 1 5634
2 2668 1 5634
2 2669 1 5634
2 2670 1 5634
2 2671 1 5655
2 2672 1 5655
2 2673 1 5655
2 2674 1 5655
2 2676 1 5655
2 2677 1 5655
2 2678 1 5655
2 2679 1 5655
2 2680 1 5655
2 2682 1 5655
2 2683 1 5655
2 2684 1 5655
2 2685 1 5655
2 2686 1 5655
2 2687 1 5655
2 2688 1 5671
2 2689 1 5671
2 2690 1 5671
2 2691 1 5671
2 2693 1 5671
2 2694 1 5671
2 2695 1 5671
2 2696 1 5671
2 2697 1 5671
2 2698 1 5671
2 2699 1 5671
2 2700 1 5671
2 2701 1 5684
2 2702 1 5684
2 2705 1 5684
2 2706 1 5684
2 2707 1 5684
2 2708 1 5692
2 2723 1 5692
2 2724 1 5692
2 2725 1 5696
2 2726 1 5696
2 2727 1 5696
2 2729 1 5700
2 2730 1 5700
2 2731 1 5703
2 2732 1 5703
2 2733 1 5703
2 2734 1 5707
2 2735 1 5707
2 2736 1 5707
2 2737 1 5711
2 2738 1 5711
2 2740 1 5736
2 2741 1 5736
2 2742 1 5739
2 2743 1 5739
2 2744 1 5742
2 2745 1 5742
2 2746 1 5745
2 2747 1 5745
2 2748 1 5756
2 2749 1 5756
2 2751 1 6025
2 2752 1 6025
2 2753 1 6028
2 2754 1 6028
2 2755 1 6031
2 2757 1 6031
2 2758 1 6034
2 2759 1 6034
2 2760 1 6037
2 2761 1 6037
2 2762 1 6040
2 2763 1 6040
2 2764 1 6045
2 2765 1 6045
2 2766 1 6048
2 2768 1 6048
2 2769 1 6051
2 2770 1 6051
2 2771 1 6054
2 2772 1 6054
2 2773 1 6080
2 2774 1 6080
2 2775 1 6091
2 2776 1 6091
2 2777 1 6108
2 2780 1 6108
2 2781 1 6117
2 2782 1 6117
2 2783 1 6140
2 2784 1 6140
2 2785 1 6149
2 2786 1 6149
2 2787 1 6164
2 2788 1 6164
2 2789 1 6168
2 2791 1 6168
2 2792 1 6175
2 2793 1 6175
2 2794 1 6197
2 2795 1 6197
2 2796 1 6200
2 2797 1 6200
2 2798 1 6203
2 2799 1 6203
2 2800 1 6206
2 2802 1 6206
2 2803 1 6209
2 2804 1 6209
2 2805 1 6212
2 2806 1 6212
2 2807 1 6215
2 2808 1 6215
2 2809 1 6218
2 2810 1 6218
2 2811 1 6238
2 2813 1 6238
2 2814 1 6241
2 2815 1 6241
2 2816 1 6244
2 2817 1 6244
2 2818 1 6247
2 2819 1 6247
2 2820 1 6250
2 2821 1 6250
2 2822 1 6253
2 2856 1 6253
2 2857 1 6256
2 2858 1 6256
2 2859 1 6259
2 2860 1 6259
2 2862 1 6262
2 2863 1 6262
2 2864 1 6265
2 2865 1 6265
2 2866 1 6268
2 2878 1 6268
2 2879 1 6271
2 2880 1 6271
2 2881 1 6274
2 2883 1 6274
2 2884 1 6277
2 2885 1 6277
2 2886 1 6280
2 2887 1 6280
2 2888 1 6283
2 2889 1 6283
2 2890 1 6286
2 2892 1 6286
2 2893 1 6289
2 2894 1 6289
2 2895 1 6292
2 2896 1 6292
2 2897 1 6295
2 2898 1 6295
2 2899 1 6298
2 2900 1 6298
2 2943 1 6301
2 2944 1 6301
2 2945 1 6304
2 2946 1 6304
2 2947 1 6307
2 2949 1 6307
2 2950 1 6310
2 2951 1 6310
2 2952 1 6313
2 2953 1 6313
2 2965 1 6316
2 2966 1 6316
2 2967 1 6319
2 2968 1 6319
2 3001 1 6322
2 3002 1 6322
2 3004 1 6325
2 3005 1 6325
2 3008 1 6328
2 3009 1 6328
2 3011 1 6331
2 3012 1 6331
2 3036 1 6335
2 3037 1 6335
2 3039 1 6338
2 3040 1 6338
2 3042 1 6341
2 3043 1 6341
2 3044 1 6344
2 3045 1 6344
2 3046 1 6347
2 3047 1 6347
2 3048 1 6350
2 3049 1 6350
2 3050 1 6353
2 3051 1 6353
2 3053 1 6356
2 3054 1 6356
2 3055 1 6359
2 3056 1 6359
2 3057 1 6364
2 3058 1 6364
2 3059 1 6367
2 3060 1 6367
2 3061 1 6370
2 3062 1 6370
2 3064 1 6397
2 3065 1 6397
2 3066 1 6411
2 3067 1 6411
2 3069 1 6415
2 3070 1 6415
2 3076 1 6415
2 3077 1 6419
2 3078 1 6419
2 3079 1 6427
2 3080 1 6427
2 3081 1 6437
2 3082 1 6437
2 3083 1 6441
2 3084 1 6441
2 3085 1 6441
2 3087 1 6445
2 3088 1 6445
2 3089 1 6466
2 3090 1 6466
2 3091 1 6478
2 3092 1 6478
2 3093 1 6482
2 3094 1 6482
2 3095 1 6486
2 3096 1 6486
2 3098 1 6490
2 3099 1 6490
2 3100 1 6494
2 3101 1 6494
2 3102 1 6500
2 3103 1 6500
2 3104 1 6504
2 3105 1 6504
2 3106 1 6508
2 3107 1 6508
2 3109 1 6512
2 3110 1 6512
2 3111 1 6516
2 3112 1 6516
2 3113 1 6526
2 3114 1 6526
2 3115 1 6536
2 3116 1 6536
2 3117 1 6539
2 3118 1 6539
2 3120 1 6553
2 3121 1 6553
2 3122 1 6556
2 3123 1 6556
2 3124 1 6566
2 3125 1 6566
2 3126 1 6569
2 3127 1 6569
2 3128 1 6572
2 3129 1 6572
2 3131 1 6575
2 3132 1 6575
2 3133 1 6580
2 3134 1 6580
2 3135 1 6584
2 3136 1 6584
2 3137 1 6587
2 3138 1 6587
2 3139 1 6592
2 3140 1 6592
2 3148 1 6599
2 3149 1 6599
2 3150 1 6606
2 3151 1 6606
2 3152 1 6609
2 3153 1 6609
2 3154 1 6619
2 3155 1 6619
2 3156 1 6622
2 3157 1 6622
2 3159 1 6634
2 3160 1 6634
2 3161 1 6637
2 3162 1 6637
2 3163 1 6724
2 3164 1 6724
2 3165 1 6792
2 3166 1 6792
2 3167 1 6795
2 3168 1 6795
2 3170 1 6817
2 3171 1 6817
2 3172 1 6817
2 3173 1 6817
2 3174 1 6817
2 3175 1 6831
2 3176 1 6831
2 3177 1 6844
2 3178 1 6844
2 3179 1 6844
2 3181 1 6844
2 3182 1 6844
2 3183 1 6857
2 3184 1 6857
2 3185 1 6866
2 3186 1 6866
2 3187 1 6866
2 3188 1 6866
2 3189 1 6866
2 3190 1 6881
2 3192 1 6881
2 3193 1 6885
2 3201 1 6885
2 3202 1 6891
2 3204 1 6891
2 3205 1 6897
2 3206 1 6897
2 3207 1 6901
2 3208 1 6901
2 3209 1 6905
2 3210 1 6905
2 3211 1 6909
2 3212 1 6909
2 3213 1 6916
2 3214 1 6916
2 3215 1 6932
2 3216 1 6932
2 3217 1 6967
2 3218 1 6967
2 3219 1 6979
2 3220 1 6979
2 3221 1 6979
2 3222 1 7003
2 3223 1 7003
2 3224 1 7006
2 3225 1 7006
2 3226 1 7023
2 3227 1 7023
2 3228 1 7023
2 3229 1 7023
2 3230 1 7028
2 3231 1 7028
2 3232 1 7031
2 3233 1 7031
2 3234 1 7034
2 3235 1 7034
2 3236 1 7037
2 3237 1 7037
2 3238 1 7041
2 3239 1 7041
2 3240 1 7049
2 3241 1 7049
2 3242 1 7049
2 3243 1 7049
2 3244 1 7054
2 3245 1 7054
2 3246 1 7057
2 3247 1 7057
2 3248 1 7060
2 3249 1 7060
2 3250 1 7065
2 3251 1 7065
2 3252 1 7076
2 3253 1 7076
2 3254 1 7080
2 3255 1 7080
2 3256 1 7090
2 3257 1 7090
2 3258 1 7094
2 3259 1 7094
2 3260 1 7097
2 3261 1 7097
2 3262 1 7101
2 3263 1 7101
2 3264 1 7190
2 3265 1 7190
2 3266 1 7190
2 3267 1 7190
2 3268 1 7190
2 3269 1 7198
2 3270 1 7198
2 3271 1 7198
2 3272 1 7198
2 3273 1 7198
2 3274 1 7209
2 3275 1 7209
2 3276 1 7212
2 3277 1 7212
2 3278 1 7219
2 3279 1 7219
2 3280 1 7222
2 3281 1 7222
2 3282 1 7225
2 3283 1 7225
2 3284 1 7236
2 3285 1 7236
2 3286 1 7239
2 3287 1 7239
2 3288 1 7242
2 3289 1 7242
2 3290 1 7245
2 3291 1 7245
2 3292 1 7250
2 3293 1 7250
2 3294 1 7250
2 3295 1 7250
2 3296 1 7250
2 3297 1 7250
2 3298 1 7257
2 3299 1 7257
2 3300 1 7260
2 3301 1 7260
2 3302 1 7263
2 3303 1 7263
2 3304 1 7270
2 3305 1 7270
2 3306 1 7270
2 3307 1 7270
2 3308 1 7270
2 3309 1 7276
2 3310 1 7276
2 3311 1 7276
2 3312 1 7276
2 3313 1 7276
2 3314 1 7282
2 3315 1 7282
2 3316 1 7282
2 3317 1 7282
2 3318 1 7282
2 3319 1 7288
2 3320 1 7288
2 3321 1 7288
2 3322 1 7288
2 3323 1 7288
2 3324 1 7294
2 3325 1 7294
2 3326 1 7294
2 3327 1 7294
2 3328 1 7294
2 3329 1 7301
2 3330 1 7301
2 3331 1 7304
2 3332 1 7304
2 3333 1 7304
2 3334 1 7304
2 3335 1 7304
2 3336 1 7310
2 3337 1 7310
2 3338 1 7310
2 3339 1 7310
2 3340 1 7310
2 3341 1 7394
2 3342 1 7394
2 3343 1 7397
2 3344 1 7397
2 3345 1 7402
2 3346 1 7402
2 3347 1 7409
2 3348 1 7409
2 3349 1 7412
2 3350 1 7412
2 3351 1 7421
2 3352 1 7421
2 3353 1 7489
2 3354 1 7489
2 3355 1 7531
2 3356 1 7531
2 3361 1 7531
2 3362 1 7531
2 3363 1 7531
2 3364 1 7537
2 3365 1 7537
2 3366 1 7537
2 3367 1 7537
2 3368 1 7537
2 3369 1 7543
2 3370 1 7543
2 3371 1 7543
2 3372 1 7543
2 3373 1 7543
2 3374 1 7549
2 3375 1 7549
2 3376 1 7549
2 3377 1 7549
2 3378 1 7549
2 3379 1 7555
2 3380 1 7555
2 3381 1 7555
2 3382 1 7555
2 3383 1 7555
2 3384 1 7561
2 3385 1 7561
2 3386 1 7561
2 3387 1 7561
2 3388 1 7561
2 3389 1 7567
2 3390 1 7567
2 3391 1 7567
2 3392 1 7567
2 3393 1 7567
2 3394 1 7573
2 3395 1 7573
2 3396 1 7573
2 3397 1 7573
2 3398 1 7573
2 3399 1 7579
2 3400 1 7579
2 3417 1 7582
2 3418 1 7582
2 3419 1 7589
2 3420 1 7589
2 3421 1 7592
2 3422 1 7592
2 3423 1 7595
2 3424 1 7595
2 3425 1 7712
2 3426 1 7712
2 3427 1 7715
2 3428 1 7715
2 3429 1 7724
2 3430 1 7724
2 3431 1 7762
2 3432 1 7762
2 3433 1 7765
2 3434 1 7765
2 3435 1 7772
2 3436 1 7772
2 3437 1 7775
2 3438 1 7775
2 3439 1 7778
2 3440 1 7778
2 3441 1 7800
2 3442 1 7800
2 3443 1 7803
2 3457 1 7803
2 3458 1 7812
2 3467 1 7812
2 3468 1 7826
2 3469 1 7826
2 3470 1 7829
2 3471 1 7829
2 3472 1 7836
2 3473 1 7836
2 3474 1 7839
2 3475 1 7839
2 3476 1 7842
2 3477 1 7842
2 3478 1 7864
2 3479 1 7864
2 3480 1 7867
2 3494 1 7867
2 3495 1 7876
2 3496 1 7876
2 3497 1 7890
2 3498 1 7890
2 3499 1 7893
2 3500 1 7893
2 3501 1 7900
2 3516 1 7900
2 3517 1 7903
2 3518 1 7903
2 3519 1 7906
2 3520 1 7906
2 3521 1 7932
2 3522 1 7932
2 3523 1 7935
2 3524 1 7935
2 3525 1 7940
2 3526 1 7940
2 3527 1 7954
2 3528 1 7954
2 3529 1 7957
2 3530 1 7957
2 3531 1 7960
2 3532 1 7960
2 3533 1 7963
2 3534 1 7963
2 3535 1 7970
2 3536 1 7970
2 3537 1 7998
2 3538 1 7998
2 3539 1 8001
2 3540 1 8001
2 3541 1 8004
2 3542 1 8004
2 3543 1 8013
2 3544 1 8013
2 3545 1 8017
2 3546 1 8017
2 3547 1 8045
2 3548 1 8045
2 3549 1 8048
2 3550 1 8048
2 3551 1 8061
2 3552 1 8061
2 3553 1 8064
2 3554 1 8064
2 3555 1 8079
2 3556 1 8079
2 3557 1 8082
2 3564 1 8082
2 3565 1 8093
2 3566 1 8093
2 3567 1 8096
2 3568 1 8096
2 3569 1 8099
2 3570 1 8099
2 3571 1 8102
2 3572 1 8102
