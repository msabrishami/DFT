1 1 0 3 0
1 5 0 3 0
1 9 0 3 0
1 13 0 3 0
1 17 0 3 0
1 21 0 3 0
1 25 0 3 0
1 29 0 3 0
1 33 0 3 0
1 37 0 3 0
1 41 0 3 0
1 45 0 3 0
1 49 0 3 0
1 53 0 3 0
1 57 0 3 0
1 61 0 3 0
1 65 0 3 0
1 69 0 3 0
1 73 0 3 0
1 77 0 3 0
1 81 0 3 0
1 85 0 3 0
1 89 0 3 0
1 93 0 3 0
1 97 0 3 0
1 101 0 3 0
1 105 0 3 0
1 109 0 3 0
1 113 0 3 0
1 117 0 3 0
1 121 0 3 0
1 125 0 3 0
1 129 0 1 0
1 130 0 1 0
1 131 0 1 0
1 132 0 1 0
1 133 0 1 0
1 134 0 1 0
1 135 0 1 0
1 136 0 1 0
1 137 0 8 0
0 250 2 1 2 2 6
0 251 2 1 2 10 14
0 252 2 1 2 18 22
0 253 2 1 2 26 30
0 254 2 1 2 34 38
0 255 2 1 2 42 46
0 256 2 1 2 50 54
0 257 2 1 2 58 62
0 258 2 1 2 66 70
0 259 2 1 2 74 78
0 260 2 1 2 82 86
0 261 2 1 2 90 94
0 262 2 1 2 98 102
0 263 2 1 2 106 110
0 264 2 1 2 114 118
0 265 2 1 2 122 126
0 266 7 1 2 129 138
0 267 7 1 2 130 139
0 268 7 1 2 131 140
0 269 7 1 2 132 141
0 270 7 1 2 133 142
0 271 7 1 2 134 143
0 272 7 1 2 135 144
0 273 7 1 2 136 145
0 274 2 1 2 3 19
0 275 2 1 2 35 51
0 276 2 1 2 7 23
0 277 2 1 2 39 55
0 278 2 1 2 11 27
0 279 2 1 2 43 59
0 280 2 1 2 15 31
0 281 2 1 2 47 63
0 282 2 1 2 67 83
0 283 2 1 2 99 115
0 284 2 1 2 71 87
0 285 2 1 2 103 119
0 286 2 1 2 75 91
0 287 2 1 2 107 123
0 288 2 1 2 79 95
0 289 2 1 2 111 127
0 290 2 2 2 250 251
0 293 2 2 2 252 253
0 296 2 2 2 254 255
0 299 2 2 2 256 257
0 302 2 2 2 258 259
0 305 2 2 2 260 261
0 308 2 2 2 262 263
0 311 2 2 2 264 265
0 314 2 1 2 274 275
0 315 2 1 2 276 277
0 316 2 1 2 278 279
0 317 2 1 2 280 281
0 318 2 1 2 282 283
0 319 2 1 2 284 285
0 320 2 1 2 286 287
0 321 2 1 2 288 289
0 338 2 1 2 146 148
0 339 2 1 2 150 152
0 340 2 1 2 147 151
0 341 2 1 2 149 153
0 342 2 1 2 154 156
0 343 2 1 2 158 160
0 344 2 1 2 155 159
0 345 2 1 2 157 161
0 346 2 1 2 266 342
0 347 2 1 2 267 343
0 348 2 1 2 268 344
0 349 2 1 2 269 345
0 350 2 1 2 270 338
0 351 2 1 2 271 339
0 352 2 1 2 272 340
0 353 2 1 2 273 341
0 354 2 12 2 314 346
0 367 2 12 2 315 347
0 380 2 12 2 316 348
0 393 2 12 2 317 349
0 406 2 12 2 318 350
0 419 2 12 2 319 351
0 432 2 12 2 320 352
0 445 2 12 2 321 353
0 554 5 1 1 162
0 555 5 1 1 174
0 556 5 1 1 186
0 557 5 1 1 163
0 558 5 1 1 175
0 559 5 1 1 198
0 560 5 1 1 164
0 561 5 1 1 187
0 562 5 1 1 199
0 563 5 1 1 176
0 564 5 1 1 188
0 565 5 1 1 200
0 566 5 1 1 222
0 567 5 1 1 246
0 568 5 1 1 223
0 569 5 1 1 234
0 570 5 1 1 210
0 571 5 1 1 247
0 572 5 1 1 211
0 573 5 1 1 235
0 574 5 1 1 212
0 575 5 1 1 224
0 576 5 1 1 236
0 577 5 1 1 213
0 578 5 1 1 225
0 579 5 1 1 248
0 580 5 1 1 214
0 581 5 1 1 237
0 582 5 1 1 249
0 583 5 1 1 226
0 584 5 1 1 238
0 585 5 1 1 291
0 586 5 1 1 177
0 587 5 1 1 201
0 588 5 1 1 178
0 589 5 1 1 189
0 590 5 1 1 165
0 591 5 1 1 202
0 592 5 1 1 166
0 593 5 1 1 190
0 594 7 1 4 554 555 556 203
0 595 7 1 4 557 558 191 559
0 596 7 1 4 560 179 561 562
0 597 7 1 4 167 563 564 565
0 598 7 1 4 574 575 576 292
0 599 7 1 4 577 578 239 579
0 600 7 1 4 580 227 581 582
0 601 7 1 4 215 583 584 585
0 602 3 4 4 594 595 596 597
0 607 3 4 4 598 599 600 601
0 620 7 4 5 216 566 240 567 303
0 625 7 4 5 217 568 569 294 304
0 630 7 4 5 570 228 241 571 306
0 635 7 4 5 572 229 573 295 307
0 640 7 4 5 168 586 192 587 309
0 645 7 4 5 169 588 589 204 310
0 650 7 4 5 590 180 193 591 312
0 655 7 4 5 592 181 593 205 313
0 692 7 1 2 170 322
0 693 7 1 2 182 323
0 694 7 1 2 194 324
0 695 7 1 2 206 325
0 696 7 1 2 171 326
0 697 7 1 2 183 327
0 698 7 1 2 195 328
0 699 7 1 2 207 329
0 700 7 1 2 172 330
0 701 7 1 2 184 331
0 702 7 1 2 196 332
0 703 7 1 2 208 333
0 704 7 1 2 173 334
0 705 7 1 2 185 335
0 706 7 1 2 197 336
0 707 7 1 2 209 337
0 708 7 1 2 218 355
0 709 7 1 2 230 356
0 710 7 1 2 242 357
0 711 7 1 2 297 358
0 712 7 1 2 219 359
0 713 7 1 2 231 360
0 714 7 1 2 243 361
0 715 7 1 2 298 362
0 716 7 1 2 220 363
0 717 7 1 2 232 364
0 718 7 1 2 244 365
0 719 7 1 2 300 366
0 720 7 1 2 221 368
0 721 7 1 2 233 369
0 722 7 1 2 245 370
0 723 7 1 2 301 371
3 724 2 0 2 4 692
3 725 2 0 2 8 693
3 726 2 0 2 12 694
3 727 2 0 2 16 695
3 728 2 0 2 20 696
3 729 2 0 2 24 697
3 730 2 0 2 28 698
3 731 2 0 2 32 699
3 732 2 0 2 36 700
3 733 2 0 2 40 701
3 734 2 0 2 44 702
3 735 2 0 2 48 703
3 736 2 0 2 52 704
3 737 2 0 2 56 705
3 738 2 0 2 60 706
3 739 2 0 2 64 707
3 740 2 0 2 68 708
3 741 2 0 2 72 709
3 742 2 0 2 76 710
3 743 2 0 2 80 711
3 744 2 0 2 84 712
3 745 2 0 2 88 713
3 746 2 0 2 92 714
3 747 2 0 2 96 715
3 748 2 0 2 100 716
3 749 2 0 2 104 717
3 750 2 0 2 108 718
3 751 2 0 2 112 719
3 752 2 0 2 116 720
3 753 2 0 2 120 721
3 754 2 0 2 124 722
3 755 2 0 2 128 723
2 2 1 1
2 3 1 1
2 4 1 1
2 6 1 5
2 7 1 5
2 8 1 5
2 10 1 9
2 11 1 9
2 12 1 9
2 14 1 13
2 15 1 13
2 16 1 13
2 18 1 17
2 19 1 17
2 20 1 17
2 22 1 21
2 23 1 21
2 24 1 21
2 26 1 25
2 27 1 25
2 28 1 25
2 30 1 29
2 31 1 29
2 32 1 29
2 34 1 33
2 35 1 33
2 36 1 33
2 38 1 37
2 39 1 37
2 40 1 37
2 42 1 41
2 43 1 41
2 44 1 41
2 46 1 45
2 47 1 45
2 48 1 45
2 50 1 49
2 51 1 49
2 52 1 49
2 54 1 53
2 55 1 53
2 56 1 53
2 58 1 57
2 59 1 57
2 60 1 57
2 62 1 61
2 63 1 61
2 64 1 61
2 66 1 65
2 67 1 65
2 68 1 65
2 70 1 69
2 71 1 69
2 72 1 69
2 74 1 73
2 75 1 73
2 76 1 73
2 78 1 77
2 79 1 77
2 80 1 77
2 82 1 81
2 83 1 81
2 84 1 81
2 86 1 85
2 87 1 85
2 88 1 85
2 90 1 89
2 91 1 89
2 92 1 89
2 94 1 93
2 95 1 93
2 96 1 93
2 98 1 97
2 99 1 97
2 100 1 97
2 102 1 101
2 103 1 101
2 104 1 101
2 106 1 105
2 107 1 105
2 108 1 105
2 110 1 109
2 111 1 109
2 112 1 109
2 114 1 113
2 115 1 113
2 116 1 113
2 118 1 117
2 119 1 117
2 120 1 117
2 122 1 121
2 123 1 121
2 124 1 121
2 126 1 125
2 127 1 125
2 128 1 125
2 138 1 137
2 139 1 137
2 140 1 137
2 141 1 137
2 142 1 137
2 143 1 137
2 144 1 137
2 145 1 137
2 146 1 290
2 147 1 290
2 148 1 293
2 149 1 293
2 150 1 296
2 151 1 296
2 152 1 299
2 153 1 299
2 154 1 302
2 155 1 302
2 156 1 305
2 157 1 305
2 158 1 308
2 159 1 308
2 160 1 311
2 161 1 311
2 162 1 354
2 163 1 354
2 164 1 354
2 165 1 354
2 166 1 354
2 167 1 354
2 168 1 354
2 169 1 354
2 170 1 354
2 171 1 354
2 172 1 354
2 173 1 354
2 174 1 367
2 175 1 367
2 176 1 367
2 177 1 367
2 178 1 367
2 179 1 367
2 180 1 367
2 181 1 367
2 182 1 367
2 183 1 367
2 184 1 367
2 185 1 367
2 186 1 380
2 187 1 380
2 188 1 380
2 189 1 380
2 190 1 380
2 191 1 380
2 192 1 380
2 193 1 380
2 194 1 380
2 195 1 380
2 196 1 380
2 197 1 380
2 198 1 393
2 199 1 393
2 200 1 393
2 201 1 393
2 202 1 393
2 203 1 393
2 204 1 393
2 205 1 393
2 206 1 393
2 207 1 393
2 208 1 393
2 209 1 393
2 210 1 406
2 211 1 406
2 212 1 406
2 213 1 406
2 214 1 406
2 215 1 406
2 216 1 406
2 217 1 406
2 218 1 406
2 219 1 406
2 220 1 406
2 221 1 406
2 222 1 419
2 223 1 419
2 224 1 419
2 225 1 419
2 226 1 419
2 227 1 419
2 228 1 419
2 229 1 419
2 230 1 419
2 231 1 419
2 232 1 419
2 233 1 419
2 234 1 432
2 235 1 432
2 236 1 432
2 237 1 432
2 238 1 432
2 239 1 432
2 240 1 432
2 241 1 432
2 242 1 432
2 243 1 432
2 244 1 432
2 245 1 432
2 246 1 445
2 247 1 445
2 248 1 445
2 249 1 445
2 291 1 445
2 292 1 445
2 294 1 445
2 295 1 445
2 297 1 445
2 298 1 445
2 300 1 445
2 301 1 445
2 303 1 602
2 304 1 602
2 306 1 602
2 307 1 602
2 309 1 607
2 310 1 607
2 312 1 607
2 313 1 607
2 322 1 620
2 323 1 620
2 324 1 620
2 325 1 620
2 326 1 625
2 327 1 625
2 328 1 625
2 329 1 625
2 330 1 630
2 331 1 630
2 332 1 630
2 333 1 630
2 334 1 635
2 335 1 635
2 336 1 635
2 337 1 635
2 355 1 640
2 356 1 640
2 357 1 640
2 358 1 640
2 359 1 645
2 360 1 645
2 361 1 645
2 362 1 645
2 363 1 650
2 364 1 650
2 365 1 650
2 366 1 650
2 368 1 655
2 369 1 655
2 370 1 655
2 371 1 655
