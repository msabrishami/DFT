1 1 0 1 0
1 2 0 2 0
2 3 1 1 2
2 4 1 2 2
1 5 0 1 0
0 6 7 2 2 1 3
2 7 1 1 6
2 8 1 1 4
2 9 1 1 4
2 10 1 1 27
2 11 1 1 27
0 12 8 2 2 7 8
2 13 1 1 12
0 14 8 2 2 11 13
2 15 1 1 14
2 16 1 1 14
0 17 5 2 1 16
2 18 1 1 28
2 19 1 1 28
2 20 1 1 17
2 21 1 1 17
0 22 5 1 1 18
0 23 8 1 2 21 9
3 24 6 0 2 10 15
3 25 3 0 2 20 22
3 26 6 0 3 23 19 5
2 27 1 2 6
2 28 1 2 12