1 0 0 7 0
1 1 0 7 0
1 2 0 7 0
1 3 0 7 0
1 4 0 7 0
1 5 0 7 0
1 6 0 7 0
1 7 0 7 0
1 8 0 7 0
1 9 0 7 0
1 10 0 7 0
1 11 0 7 0
1 12 0 7 0
1 13 0 7 0
1 14 0 7 0
1 15 0 7 0
1 16 0 7 0
1 17 0 7 0
1 18 0 7 0
1 19 0 7 0
1 20 0 7 0
1 21 0 7 0
1 22 0 7 0
1 23 0 7 0
1 24 0 7 0
1 25 0 7 0
1 26 0 7 0
1 27 0 7 0
1 28 0 7 0
1 29 0 7 0
1 30 0 7 0
1 31 0 7 0
1 32 0 3 0
1 33 0 3 0
1 34 0 3 0
1 35 0 3 0
1 36 0 3 0
1 37 0 3 0
1 38 0 3 0
1 39 0 2 0
1 40 0 17 0
2 41 1 0 
2 42 1 0 
2 43 1 0 
2 44 1 0 
2 45 1 0 
2 46 1 0 
2 47 1 0 
2 48 1 1 
2 49 1 1 
2 50 1 1 
2 51 1 1 
2 52 1 1 
2 53 1 1 
2 54 1 1 
2 55 1 2 
2 56 1 2 
2 57 1 2 
2 58 1 2 
2 59 1 2 
2 60 1 2 
2 61 1 2 
2 62 1 3 
2 63 1 3 
2 64 1 3 
2 65 1 3 
2 66 1 3 
2 67 1 3 
2 68 1 3 
2 69 1 4 
2 70 1 4 
2 71 1 4 
2 72 1 4 
2 73 1 4 
2 74 1 4 
2 75 1 4 
2 76 1 5 
2 77 1 5 
2 78 1 5 
2 79 1 5 
2 80 1 5 
2 81 1 5 
2 82 1 5 
2 83 1 6 
2 84 1 6 
2 85 1 6 
2 86 1 6 
2 87 1 6 
2 88 1 6 
2 89 1 6 
2 90 1 7 
2 91 1 7 
2 92 1 7 
2 93 1 7 
2 94 1 7 
2 95 1 7 
2 96 1 7 
2 97 1 8 
2 98 1 8 
2 99 1 8 
2 100 1 8 
2 101 1 8 
2 102 1 8 
2 103 1 8 
2 104 1 9 
2 105 1 9 
2 106 1 9 
2 107 1 9 
2 108 1 9 
2 109 1 9 
2 110 1 9 
2 111 1 10 
2 112 1 10 
2 113 1 10 
2 114 1 10 
2 115 1 10 
2 116 1 10 
2 117 1 10 
2 118 1 11 
2 119 1 11 
2 120 1 11 
2 121 1 11 
2 122 1 11 
2 123 1 11 
2 124 1 11 
2 125 1 12 
2 126 1 12 
2 127 1 12 
2 128 1 12 
2 129 1 12 
2 130 1 12 
2 131 1 12 
2 132 1 13 
2 133 1 13 
2 134 1 13 
2 135 1 13 
2 136 1 13 
2 137 1 13 
2 138 1 13 
2 139 1 14 
2 140 1 14 
2 141 1 14 
2 142 1 14 
2 143 1 14 
2 144 1 14 
2 145 1 14 
2 146 1 15 
2 147 1 15 
2 148 1 15 
2 149 1 15 
2 150 1 15 
2 151 1 15 
2 152 1 15 
2 153 1 16 
2 154 1 16 
2 155 1 16 
2 156 1 16 
2 157 1 16 
2 158 1 16 
2 159 1 16 
2 160 1 17 
2 161 1 17 
2 162 1 17 
2 163 1 17 
2 164 1 17 
2 165 1 17 
2 166 1 17 
2 167 1 18 
2 168 1 18 
2 169 1 18 
2 170 1 18 
2 171 1 18 
2 172 1 18 
2 173 1 18 
2 174 1 19 
2 175 1 19 
2 176 1 19 
2 177 1 19 
2 178 1 19 
2 179 1 19 
2 180 1 19 
2 181 1 20 
2 182 1 20 
2 183 1 20 
2 184 1 20 
2 185 1 20 
2 186 1 20 
2 187 1 20 
2 188 1 21 
2 189 1 21 
2 190 1 21 
2 191 1 21 
2 192 1 21 
2 193 1 21 
2 194 1 21 
2 195 1 22 
2 196 1 22 
2 197 1 22 
2 198 1 22 
2 199 1 22 
2 200 1 22 
2 201 1 22 
2 202 1 23 
2 203 1 23 
2 204 1 23 
2 205 1 23 
2 206 1 23 
2 207 1 23 
2 208 1 23 
2 209 1 24 
2 210 1 24 
2 211 1 24 
2 212 1 24 
2 213 1 24 
2 214 1 24 
2 215 1 24 
2 216 1 25 
2 217 1 25 
2 218 1 25 
2 219 1 25 
2 220 1 25 
2 221 1 25 
2 222 1 25 
2 223 1 26 
2 224 1 26 
2 225 1 26 
2 226 1 26 
2 227 1 26 
2 228 1 26 
2 229 1 26 
2 230 1 27 
2 231 1 27 
2 232 1 27 
2 233 1 27 
2 234 1 27 
2 235 1 27 
2 236 1 27 
2 237 1 28 
2 238 1 28 
2 239 1 28 
2 240 1 28 
2 241 1 28 
2 242 1 28 
2 243 1 28 
2 244 1 29 
2 245 1 29 
2 246 1 29 
2 247 1 29 
2 248 1 29 
2 249 1 29 
2 250 1 29 
2 251 1 30 
2 252 1 30 
2 253 1 30 
2 254 1 30 
2 255 1 30 
2 256 1 30 
2 257 1 30 
2 258 1 31 
2 259 1 31 
2 260 1 31 
2 261 1 31 
2 262 1 31 
2 263 1 31 
2 264 1 31 
2 265 1 32 
2 266 1 32 
2 267 1 32 
2 268 1 33 
2 269 1 33 
2 270 1 33 
2 271 1 34 
2 272 1 34 
2 273 1 34 
2 274 1 35 
2 275 1 35 
2 276 1 35 
2 277 1 36 
2 278 1 36 
2 279 1 36 
2 280 1 37 
2 281 1 37 
2 282 1 37 
2 283 1 38 
2 284 1 38 
2 285 1 38 
2 286 1 39 
2 287 1 39 
2 288 1 40 
2 289 1 40 
2 290 1 40 
2 291 1 40 
2 292 1 40 
2 293 1 40 
2 294 1 40 
2 295 1 40 
2 296 1 40 
2 297 1 40 
2 298 1 40 
2 299 1 40 
2 300 1 40 
2 301 1 40 
2 302 1 40 
2 303 1 40 
2 304 1 40 
0 305 5 2 1 286
0 306 6 1 2 287 289
0 307 7 1 2 280 290
0 308 6 1 2 282 291
0 309 7 1 2 274 292
0 310 6 1 2 276 293
0 311 5 4 1 151
0 312 7 1 2 271 294
0 313 6 1 2 273 295
0 314 5 4 1 145
0 315 7 1 2 268 296
0 316 6 1 2 270 297
0 317 5 4 1 250
0 318 5 4 1 264
0 319 5 4 1 236
0 320 5 4 1 222
0 321 5 4 1 138
0 322 7 1 2 265 298
0 323 6 1 2 267 299
0 324 5 4 1 166
0 325 5 4 1 180
0 326 5 4 1 194
0 327 5 4 1 208
0 328 5 4 1 131
0 329 7 1 2 277 300
0 330 6 1 2 279 301
0 331 5 4 1 74
0 332 5 4 1 82
0 333 5 4 1 88
0 334 5 4 1 96
0 335 5 4 1 158
0 336 5 4 1 187
0 337 5 4 1 214
0 338 5 4 1 243
0 339 7 1 2 283 302
0 340 5 8 1 303
0 341 6 1 2 285 304
0 342 5 4 1 46
0 343 5 4 1 61
0 344 5 4 1 67
0 345 5 4 1 54
0 346 5 4 1 116
0 347 5 4 1 124
0 348 5 4 1 102
0 349 5 4 1 110
0 350 5 4 1 172
0 351 5 4 1 201
0 352 5 4 1 228
0 353 5 4 1 257
2 354 1 305 
2 355 1 305 
2 356 1 311 
2 357 1 311 
2 358 1 311 
2 359 1 311 
2 360 1 314 
2 361 1 314 
2 362 1 314 
2 363 1 314 
2 364 1 317 
2 365 1 317 
2 366 1 317 
2 367 1 317 
2 368 1 318 
2 369 1 318 
2 370 1 318 
2 371 1 318 
2 372 1 319 
2 373 1 319 
2 374 1 319 
2 375 1 319 
2 376 1 320 
2 377 1 320 
2 378 1 320 
2 379 1 320 
2 380 1 321 
2 381 1 321 
2 382 1 321 
2 383 1 321 
2 384 1 324 
2 385 1 324 
2 386 1 324 
2 387 1 324 
2 388 1 325 
2 389 1 325 
2 390 1 325 
2 391 1 325 
2 392 1 326 
2 393 1 326 
2 394 1 326 
2 395 1 326 
2 396 1 327 
2 397 1 327 
2 398 1 327 
2 399 1 327 
2 400 1 328 
2 401 1 328 
2 402 1 328 
2 403 1 328 
2 404 1 331 
2 405 1 331 
2 406 1 331 
2 407 1 331 
2 408 1 332 
2 409 1 332 
2 410 1 332 
2 411 1 332 
2 412 1 333 
2 413 1 333 
2 414 1 333 
2 415 1 333 
2 416 1 334 
2 417 1 334 
2 418 1 334 
2 419 1 334 
2 420 1 335 
2 421 1 335 
2 422 1 335 
2 423 1 335 
2 424 1 336 
2 425 1 336 
2 426 1 336 
2 427 1 336 
2 428 1 337 
2 429 1 337 
2 430 1 337 
2 431 1 337 
2 432 1 338 
2 433 1 338 
2 434 1 338 
2 435 1 338 
2 436 1 340 
2 437 1 340 
2 438 1 340 
2 439 1 340 
2 440 1 340 
2 441 1 340 
2 442 1 340 
2 443 1 340 
2 444 1 342 
2 445 1 342 
2 446 1 342 
2 447 1 342 
2 448 1 343 
2 449 1 343 
2 450 1 343 
2 451 1 343 
2 452 1 344 
2 453 1 344 
2 454 1 344 
2 455 1 344 
2 456 1 345 
2 457 1 345 
2 458 1 345 
2 459 1 345 
2 460 1 346 
2 461 1 346 
2 462 1 346 
2 463 1 346 
2 464 1 347 
2 465 1 347 
2 466 1 347 
2 467 1 347 
2 468 1 348 
2 469 1 348 
2 470 1 348 
2 471 1 348 
2 472 1 349 
2 473 1 349 
2 474 1 349 
2 475 1 349 
2 476 1 350 
2 477 1 350 
2 478 1 350 
2 479 1 350 
2 480 1 351 
2 481 1 351 
2 482 1 351 
2 483 1 351 
2 484 1 352 
2 485 1 352 
2 486 1 352 
2 487 1 352 
2 488 1 353 
2 489 1 353 
2 490 1 353 
2 491 1 353 
0 492 4 1 2 354 436
0 493 6 1 2 260 372
0 494 6 1 2 232 368
0 495 4 1 2 204 388
0 496 4 1 2 176 396
0 497 6 1 2 205 389
0 498 6 1 2 177 397
0 499 4 1 2 261 373
0 500 4 1 2 233 369
0 501 6 1 2 141 380
0 502 6 1 2 134 360
0 503 4 1 2 127 356
0 504 4 1 2 148 400
0 505 6 1 2 128 357
0 506 6 1 2 149 401
0 507 4 1 2 142 381
0 508 4 1 2 135 361
0 509 6 1 2 246 376
0 510 6 1 2 218 364
0 511 4 1 2 190 384
0 512 4 1 2 162 392
0 513 6 1 2 191 385
0 514 6 1 2 163 393
0 515 4 1 2 247 377
0 516 4 1 2 219 365
0 517 6 1 2 120 416
0 518 6 1 2 92 464
0 519 4 1 2 64 358
0 520 4 1 2 150 452
0 521 6 1 2 65 359
0 522 6 1 2 152 453
0 523 4 1 2 121 417
0 524 4 1 2 93 465
0 525 6 1 2 143 460
0 526 6 1 2 113 362
0 527 4 1 2 85 448
0 528 4 1 2 57 412
0 529 6 1 2 86 449
0 530 6 1 2 58 413
0 531 4 1 2 144 461
0 532 4 1 2 114 363
0 533 6 1 2 262 488
0 534 6 1 2 253 370
0 535 4 1 2 248 432
0 536 4 1 2 239 366
0 537 6 1 2 249 433
0 538 6 1 2 240 367
0 539 4 1 2 263 489
0 540 4 1 2 254 371
0 541 6 1 2 220 428
0 542 6 1 2 211 378
0 543 4 1 2 234 484
0 544 4 1 2 225 374
0 545 6 1 2 235 485
0 546 6 1 2 226 375
0 547 4 1 2 221 429
0 548 4 1 2 212 379
0 549 6 1 2 136 456
0 550 6 1 2 50 382
0 551 4 1 2 106 408
0 552 4 1 2 78 472
0 553 6 1 2 107 409
0 554 6 1 2 79 473
0 555 4 1 2 137 457
0 556 4 1 2 51 383
0 557 6 1 2 178 476
0 558 6 1 2 169 390
0 559 4 1 2 164 420
0 560 4 1 2 155 386
0 561 6 1 2 165 421
0 562 6 1 2 156 387
0 563 4 1 2 179 477
0 564 4 1 2 170 391
0 565 6 1 2 206 480
0 566 6 1 2 197 398
0 567 4 1 2 192 424
0 568 4 1 2 183 394
0 569 6 1 2 193 425
0 570 6 1 2 184 395
0 571 4 1 2 207 481
0 572 4 1 2 198 399
0 573 6 1 2 129 468
0 574 6 1 2 99 402
0 575 4 1 2 71 444
0 576 4 1 2 43 404
0 577 6 1 2 72 445
0 578 6 1 2 44 405
0 579 4 1 2 130 469
0 580 4 1 2 100 403
0 581 6 1 2 94 414
0 582 6 1 2 87 418
0 583 4 1 2 80 406
0 584 4 1 2 73 410
0 585 6 1 2 81 407
0 586 6 1 2 75 411
0 587 4 1 2 95 415
0 588 4 1 2 89 419
0 589 6 1 2 241 430
0 590 6 1 2 213 434
0 591 4 1 2 185 422
0 592 4 1 2 157 426
0 593 6 1 2 186 423
0 594 6 1 2 159 427
0 595 4 1 2 242 431
0 596 4 1 2 215 435
0 597 6 1 2 52 454
0 598 6 1 2 66 458
0 599 4 1 2 59 446
0 600 4 1 2 45 450
0 601 6 1 2 60 447
0 602 6 1 2 47 451
0 603 4 1 2 53 455
0 604 4 1 2 68 459
0 605 6 1 2 108 470
0 606 6 1 2 101 474
0 607 4 1 2 122 462
0 608 4 1 2 115 466
0 609 6 1 2 123 463
0 610 6 1 2 117 467
0 611 4 1 2 109 471
0 612 4 1 2 103 475
0 613 6 1 2 255 486
0 614 6 1 2 227 490
0 615 4 1 2 199 478
0 616 4 1 2 171 482
0 617 6 1 2 200 479
0 618 6 1 2 173 483
0 619 4 1 2 256 487
0 620 4 1 2 229 491
0 621 6 1 2 494 493
0 622 4 1 2 496 495
0 623 6 1 2 498 497
0 624 4 1 2 500 499
0 625 6 1 2 502 501
0 626 4 1 2 504 503
0 627 6 1 2 506 505
0 628 4 1 2 508 507
0 629 6 1 2 510 509
0 630 4 1 2 512 511
0 631 6 1 2 514 513
0 632 4 1 2 516 515
0 633 6 1 2 518 517
0 634 4 1 2 520 519
0 635 6 1 2 522 521
0 636 4 1 2 524 523
0 637 6 1 2 526 525
0 638 4 1 2 528 527
0 639 6 1 2 530 529
0 640 4 1 2 532 531
0 641 6 1 2 534 533
0 642 4 1 2 536 535
0 643 6 1 2 538 537
0 644 4 1 2 540 539
0 645 6 1 2 542 541
0 646 4 1 2 544 543
0 647 6 1 2 546 545
0 648 4 1 2 548 547
0 649 6 1 2 550 549
0 650 4 1 2 552 551
0 651 6 1 2 554 553
0 652 4 1 2 556 555
0 653 6 1 2 558 557
0 654 4 1 2 560 559
0 655 6 1 2 562 561
0 656 4 1 2 564 563
0 657 6 1 2 566 565
0 658 4 1 2 568 567
0 659 6 1 2 570 569
0 660 4 1 2 572 571
0 661 6 1 2 574 573
0 662 4 1 2 576 575
0 663 6 1 2 578 577
0 664 4 1 2 580 579
0 665 6 1 2 582 581
0 666 4 1 2 584 583
0 667 6 1 2 586 585
0 668 4 1 2 588 587
0 669 6 1 2 590 589
0 670 4 1 2 592 591
0 671 6 1 2 594 593
0 672 4 1 2 596 595
0 673 6 1 2 598 597
0 674 4 1 2 600 599
0 675 6 1 2 602 601
0 676 4 1 2 604 603
0 677 6 1 2 606 605
0 678 4 1 2 608 607
0 679 6 1 2 610 609
0 680 4 1 2 612 611
0 681 6 1 2 614 613
0 682 4 1 2 616 615
0 683 6 1 2 618 617
0 684 4 1 2 620 619
0 685 6 2 2 622 621
0 686 6 2 2 624 623
0 687 6 1 2 626 625
0 688 6 1 2 628 627
0 689 6 2 2 630 629
0 690 6 2 2 632 631
0 691 6 2 2 634 633
0 692 6 2 2 636 635
0 693 6 2 2 638 637
0 694 6 2 2 640 639
0 695 6 1 2 642 641
0 696 6 1 2 644 643
0 697 6 1 2 646 645
0 698 6 1 2 648 647
0 699 6 2 2 650 649
0 700 6 2 2 652 651
0 701 6 1 2 654 653
0 702 6 1 2 656 655
0 703 6 1 2 658 657
0 704 6 1 2 660 659
0 705 6 2 2 662 661
0 706 6 2 2 664 663
0 707 6 1 2 666 665
0 708 6 1 2 668 667
0 709 6 2 2 670 669
0 710 6 2 2 672 671
0 711 6 1 2 674 673
0 712 6 1 2 676 675
0 713 6 1 2 678 677
0 714 6 1 2 680 679
0 715 6 2 2 682 681
0 716 6 2 2 684 683
0 717 6 3 2 688 687
0 718 6 3 2 696 695
0 719 6 3 2 698 697
0 720 6 3 2 702 701
0 721 6 3 2 704 703
0 722 6 3 2 708 707
0 723 6 3 2 712 711
0 724 6 3 2 714 713
2 725 1 685 
2 726 1 685 
2 727 1 686 
2 728 1 686 
2 729 1 689 
2 730 1 689 
2 731 1 690 
2 732 1 690 
2 733 1 691 
2 734 1 691 
2 735 1 692 
2 736 1 692 
2 737 1 693 
2 738 1 693 
2 739 1 694 
2 740 1 694 
2 741 1 699 
2 742 1 699 
2 743 1 700 
2 744 1 700 
2 745 1 705 
2 746 1 705 
2 747 1 706 
2 748 1 706 
2 749 1 709 
2 750 1 709 
2 751 1 710 
2 752 1 710 
2 753 1 715 
2 754 1 715 
2 755 1 716 
2 756 1 716 
0 757 6 1 2 725 727
0 758 7 1 2 726 728
0 759 6 1 2 729 731
0 760 7 1 2 730 732
0 761 6 1 2 733 735
0 762 7 1 2 734 736
0 763 6 1 2 737 739
0 764 7 1 2 738 740
0 765 6 1 2 741 743
0 766 7 1 2 742 744
0 767 6 1 2 745 747
0 768 7 1 2 746 748
0 769 6 1 2 749 751
0 770 7 1 2 750 752
0 771 6 1 2 753 755
0 772 7 1 2 754 756
2 773 1 717 
2 774 1 717 
2 775 1 717 
2 776 1 718 
2 777 1 718 
2 778 1 718 
2 779 1 719 
2 780 1 719 
2 781 1 719 
2 782 1 720 
2 783 1 720 
2 784 1 720 
2 785 1 721 
2 786 1 721 
2 787 1 721 
2 788 1 722 
2 789 1 722 
2 790 1 722 
2 791 1 723 
2 792 1 723 
2 793 1 723 
2 794 1 724 
2 795 1 724 
2 796 1 724 
0 797 5 2 1 774
0 798 5 2 1 777
0 799 5 2 1 781
0 800 5 2 1 783
0 801 5 2 1 787
0 802 5 2 1 789
0 803 5 2 1 792
0 804 5 2 1 796
2 805 1 797 
2 806 1 797 
2 807 1 798 
2 808 1 798 
2 809 1 799 
2 810 1 799 
2 811 1 800 
2 812 1 800 
2 813 1 801 
2 814 1 801 
2 815 1 802 
2 816 1 802 
2 817 1 803 
2 818 1 803 
2 819 1 804 
2 820 1 804 
0 821 6 1 2 773 815
0 822 6 1 2 805 788
0 823 6 1 2 806 794
0 824 6 1 2 775 819
0 825 6 1 2 776 813
0 826 6 1 2 807 785
0 827 6 1 2 779 811
0 828 6 1 2 809 782
0 829 6 1 2 808 780
0 830 6 1 2 778 810
0 831 6 1 2 812 786
0 832 6 1 2 784 814
0 833 6 1 2 816 791
0 834 6 1 2 790 817
0 835 6 1 2 818 795
0 836 6 1 2 793 820
0 837 6 2 2 822 821
0 838 6 2 2 824 823
0 839 6 2 2 826 825
0 840 6 2 2 828 827
0 841 6 2 2 830 829
0 842 6 2 2 832 831
0 843 6 2 2 834 833
0 844 6 2 2 836 835
2 845 1 837 
2 846 1 837 
2 847 1 838 
2 848 1 838 
2 849 1 839 
2 850 1 839 
2 851 1 840 
2 852 1 840 
2 853 1 841 
2 854 1 841 
2 855 1 842 
2 856 1 842 
2 857 1 843 
2 858 1 843 
2 859 1 844 
2 860 1 844 
0 861 4 1 2 492 845
0 862 5 2 1 846
0 863 4 1 2 307 847
0 864 5 2 1 848
0 865 4 1 2 309 849
0 866 5 2 1 850
0 867 4 1 2 312 851
0 868 5 2 1 852
0 869 4 1 2 315 853
0 870 5 2 1 854
0 871 4 1 2 322 855
0 872 5 2 1 856
0 873 4 1 2 329 857
0 874 5 2 1 858
0 875 4 1 2 339 859
0 876 5 2 1 860
2 877 1 862 
2 878 1 862 
2 879 1 864 
2 880 1 864 
2 881 1 866 
2 882 1 866 
2 883 1 868 
2 884 1 868 
2 885 1 870 
2 886 1 870 
2 887 1 872 
2 888 1 872 
2 889 1 874 
2 890 1 874 
2 891 1 876 
2 892 1 876 
0 893 4 1 2 355 877
0 894 6 1 2 306 878
0 895 4 1 2 879 437
0 896 6 1 2 308 880
0 897 4 1 2 881 438
0 898 6 1 2 310 882
0 899 4 1 2 883 439
0 900 6 1 2 313 884
0 901 4 1 2 885 440
0 902 6 1 2 316 886
0 903 4 1 2 887 441
0 904 6 1 2 323 888
0 905 4 1 2 889 442
0 906 6 1 2 330 890
0 907 4 1 2 443 891
0 908 6 1 2 341 892
0 909 6 2 2 893 288
0 910 6 2 2 895 281
0 911 6 2 2 897 275
0 912 6 2 2 899 272
0 913 6 2 2 901 269
0 914 6 2 2 903 266
0 915 6 2 2 905 278
0 916 6 2 2 907 284
2 917 1 909 
2 918 1 909 
2 919 1 910 
2 920 1 910 
2 921 1 911 
2 922 1 911 
2 923 1 912 
2 924 1 912 
2 925 1 913 
2 926 1 913 
2 927 1 914 
2 928 1 914 
2 929 1 915 
2 930 1 915 
2 931 1 916 
2 932 1 916 
0 933 5 1 1 917
0 934 6 1 2 894 918
0 935 5 1 1 919
0 936 6 1 2 896 920
0 937 5 1 1 921
0 938 6 1 2 898 922
0 939 5 1 1 923
0 940 6 1 2 900 924
0 941 5 1 1 925
0 942 6 1 2 902 926
0 943 5 1 1 927
0 944 6 1 2 904 928
0 945 5 1 1 929
0 946 6 1 2 906 930
0 947 5 1 1 931
0 948 6 1 2 908 932
0 949 4 1 2 933 861
0 950 6 1 2 758 934
0 951 4 1 2 935 863
0 952 6 1 2 760 936
0 953 4 1 2 937 865
0 954 6 1 2 762 938
0 955 4 1 2 939 867
0 956 6 1 2 764 940
0 957 4 1 2 941 869
0 958 6 1 2 766 942
0 959 4 1 2 943 871
0 960 6 1 2 768 944
0 961 4 1 2 945 873
0 962 6 1 2 770 946
0 963 4 1 2 947 875
0 964 6 1 2 772 948
0 965 6 1 2 949 757
0 966 6 1 2 951 759
0 967 6 1 2 953 761
0 968 6 1 2 955 763
0 969 6 1 2 957 765
0 970 6 1 2 959 767
0 971 6 1 2 961 769
0 972 6 1 2 963 771
0 973 6 3 2 950 965
0 974 6 4 2 952 966
0 975 6 5 2 954 967
0 976 6 2 2 956 968
0 977 6 2 2 958 969
0 978 6 3 2 960 970
0 979 6 4 2 962 971
0 980 6 5 2 964 972
2 981 1 973 
2 982 1 973 
2 983 1 973 
2 984 1 974 
2 985 1 974 
2 986 1 974 
2 987 1 974 
2 988 1 975 
2 989 1 975 
2 990 1 975 
2 991 1 975 
2 992 1 975 
2 993 1 976 
2 994 1 976 
2 995 1 977 
2 996 1 977 
2 997 1 978 
2 998 1 978 
2 999 1 978 
2 1000 1 979 
2 1001 1 979 
2 1002 1 979 
2 1003 1 979 
2 1004 1 980 
2 1005 1 980 
2 1006 1 980 
2 1007 1 980 
2 1008 1 980 
0 1009 6 1 2 993 997
0 1010 4 1 2 988 995
0 1011 5 6 1 1000
0 1012 6 1 2 981 1001
0 1013 4 1 2 985 1006
0 1014 5 6 1 982
0 1015 5 5 1 1007
0 1016 5 6 1 986
0 1017 5 5 1 990
0 1018 6 2 2 983 987
0 1019 5 7 1 994
0 1020 5 8 1 996
0 1021 5 7 1 999
0 1022 4 1 2 1003 1008
2 1023 1 1011 
2 1024 1 1011 
2 1025 1 1011 
2 1026 1 1011 
2 1027 1 1011 
2 1028 1 1011 
2 1029 1 1014 
2 1030 1 1014 
2 1031 1 1014 
2 1032 1 1014 
2 1033 1 1014 
2 1034 1 1014 
2 1035 1 1015 
2 1036 1 1015 
2 1037 1 1015 
2 1038 1 1015 
2 1039 1 1015 
2 1040 1 1016 
2 1041 1 1016 
2 1042 1 1016 
2 1043 1 1016 
2 1044 1 1016 
2 1045 1 1016 
2 1046 1 1017 
2 1047 1 1017 
2 1048 1 1017 
2 1049 1 1017 
2 1050 1 1017 
2 1051 1 1018 
2 1052 1 1018 
2 1053 1 1019 
2 1054 1 1019 
2 1055 1 1019 
2 1056 1 1019 
2 1057 1 1019 
2 1058 1 1019 
2 1059 1 1019 
2 1060 1 1020 
2 1061 1 1020 
2 1062 1 1020 
2 1063 1 1020 
2 1064 1 1020 
2 1065 1 1020 
2 1066 1 1020 
2 1067 1 1020 
2 1068 1 1021 
2 1069 1 1021 
2 1070 1 1021 
2 1071 1 1021 
2 1072 1 1021 
2 1073 1 1021 
2 1074 1 1021 
0 1075 6 1 2 1060 998
0 1076 6 1 2 1033 1044
0 1077 5 2 1 1051
0 1078 4 1 2 1028 984
0 1079 4 1 2 1045 1002
0 1080 6 1 2 1058 1066
0 1081 4 3 2 1059 1067
2 1082 1 1077 
2 1083 1 1077 
2 1084 1 1081 
2 1085 1 1081 
2 1086 1 1081 
0 1087 7 1 2 1084 1068
0 1088 6 1 2 1082 1004
0 1089 4 1 2 1083 1005
0 1090 6 1 2 991 1085
0 1091 4 1 2 992 1086
0 1092 4 1 2 1089 1027
0 1093 4 1 2 1091 1074
0 1094 6 1 2 1092 1076
0 1095 6 1 2 1093 1080
0 1096 7 3 2 1094 1088
0 1097 7 3 2 1095 1090
2 1098 1 1096 
2 1099 1 1096 
2 1100 1 1096 
2 1101 1 1097 
2 1102 1 1097 
2 1103 1 1097 
0 1104 4 1 2 1009 1098
0 1105 4 1 2 1099 989
0 1106 4 1 2 1100 1046
0 1107 4 1 2 1012 1101
0 1108 4 1 2 1039 1102
0 1109 4 1 2 1052 1103
0 1110 7 4 2 1010 1104
0 1111 7 4 2 1087 1105
0 1112 6 2 2 1106 1053
0 1113 7 4 2 1013 1107
0 1114 7 2 2 1108 1034
0 1115 7 4 2 1022 1109
2 1116 1 1110 
2 1117 1 1110 
2 1118 1 1110 
2 1119 1 1110 
2 1120 1 1111 
2 1121 1 1111 
2 1122 1 1111 
2 1123 1 1111 
2 1124 1 1112 
2 1125 1 1112 
2 1126 1 1113 
2 1127 1 1113 
2 1128 1 1113 
2 1129 1 1113 
2 1130 1 1114 
2 1131 1 1114 
2 1132 1 1115 
2 1133 1 1115 
2 1134 1 1115 
2 1135 1 1115 
0 1136 6 2 2 1116 1029
0 1137 6 2 2 1117 1035
0 1138 6 2 2 1118 1040
0 1139 6 2 2 1119 1023
0 1140 4 4 2 1075 1124
0 1141 6 2 2 1120 1031
0 1142 6 2 2 1121 1037
0 1143 6 2 2 1122 1042
0 1144 6 2 2 1123 1025
0 1145 4 1 2 1125 1061
0 1146 7 4 2 1078 1130
0 1147 6 2 2 1126 1048
0 1148 6 2 2 1127 1055
0 1149 6 2 2 1128 1063
0 1150 6 2 2 1129 1071
0 1151 7 4 2 1079 1131
0 1152 6 2 2 1050 1132
0 1153 6 2 2 1133 1057
0 1154 6 2 2 1134 1065
0 1155 6 2 2 1135 1073
0 1156 7 4 2 1145 1069
2 1157 1 1136 
2 1158 1 1136 
2 1159 1 1137 
2 1160 1 1137 
2 1161 1 1138 
2 1162 1 1138 
2 1163 1 1139 
2 1164 1 1139 
2 1165 1 1140 
2 1166 1 1140 
2 1167 1 1140 
2 1168 1 1140 
2 1169 1 1141 
2 1170 1 1141 
2 1171 1 1142 
2 1172 1 1142 
2 1173 1 1143 
2 1174 1 1143 
2 1175 1 1144 
2 1176 1 1144 
2 1177 1 1146 
2 1178 1 1146 
2 1179 1 1146 
2 1180 1 1146 
2 1181 1 1147 
2 1182 1 1147 
2 1183 1 1148 
2 1184 1 1148 
2 1185 1 1149 
2 1186 1 1149 
2 1187 1 1150 
2 1188 1 1150 
2 1189 1 1151 
2 1190 1 1151 
2 1191 1 1151 
2 1192 1 1151 
2 1193 1 1152 
2 1194 1 1152 
2 1195 1 1153 
2 1196 1 1153 
2 1197 1 1154 
2 1198 1 1154 
2 1199 1 1155 
2 1200 1 1155 
0 1201 6 1 2 258 1157
0 1202 3 1 2 259 1158
0 1203 6 1 2 251 1159
0 1204 3 1 2 252 1160
0 1205 6 1 2 244 1161
0 1206 3 1 2 245 1162
0 1207 6 1 2 237 1163
0 1208 3 1 2 238 1164
0 1209 6 2 2 1165 1030
0 1210 6 2 2 1166 1036
0 1211 6 2 2 1167 1041
0 1212 6 2 2 1168 1024
0 1213 6 1 2 202 1169
0 1214 3 1 2 203 1170
0 1215 6 1 2 195 1171
0 1216 3 1 2 196 1172
0 1217 6 1 2 188 1173
0 1218 3 1 2 189 1174
0 1219 6 1 2 181 1175
0 1220 3 1 2 182 1176
0 1221 6 2 2 1177 1047
0 1222 6 2 2 1178 1054
0 1223 6 2 2 1179 1062
0 1224 6 2 2 1180 1070
0 1225 6 1 2 118 1181
0 1226 3 1 2 119 1182
0 1227 6 1 2 111 1183
0 1228 3 1 2 112 1184
0 1229 6 1 2 104 1185
0 1230 3 1 2 105 1186
0 1231 6 1 2 97 1187
0 1232 3 1 2 98 1188
0 1233 6 2 2 1189 1049
0 1234 6 2 2 1190 1056
0 1235 6 2 2 1191 1064
0 1236 6 2 2 1192 1072
0 1237 6 1 2 62 1193
0 1238 3 1 2 63 1194
0 1239 6 1 2 55 1195
0 1240 3 1 2 56 1196
0 1241 6 1 2 48 1197
0 1242 3 1 2 49 1198
0 1243 6 1 2 41 1199
0 1244 3 1 2 42 1200
2 1245 1 1156 
2 1246 1 1156 
2 1247 1 1156 
2 1248 1 1156 
3 1249 6 0 2 1202 1201
3 1250 6 0 2 1204 1203
3 1251 6 0 2 1206 1205
3 1252 6 0 2 1208 1207
3 1253 6 0 2 1214 1213
3 1254 6 0 2 1216 1215
3 1255 6 0 2 1218 1217
3 1256 6 0 2 1220 1219
0 1257 6 2 2 1245 1032
0 1258 6 2 2 1246 1038
0 1259 6 2 2 1247 1043
0 1260 6 2 2 1248 1026
3 1261 6 0 2 1226 1225
3 1262 6 0 2 1228 1227
3 1263 6 0 2 1230 1229
3 1264 6 0 2 1232 1231
3 1265 6 0 2 1238 1237
3 1266 6 0 2 1240 1239
3 1267 6 0 2 1242 1241
3 1268 6 0 2 1244 1243
2 1269 1 1209 
2 1270 1 1209 
2 1271 1 1210 
2 1272 1 1210 
2 1273 1 1211 
2 1274 1 1211 
2 1275 1 1212 
2 1276 1 1212 
2 1277 1 1221 
2 1278 1 1221 
2 1279 1 1222 
2 1280 1 1222 
2 1281 1 1223 
2 1282 1 1223 
2 1283 1 1224 
2 1284 1 1224 
2 1285 1 1233 
2 1286 1 1233 
2 1287 1 1234 
2 1288 1 1234 
2 1289 1 1235 
2 1290 1 1235 
2 1291 1 1236 
2 1292 1 1236 
0 1293 6 1 2 230 1269
0 1294 3 1 2 231 1270
0 1295 6 1 2 223 1271
0 1296 3 1 2 224 1272
0 1297 6 1 2 216 1273
0 1298 3 1 2 217 1274
0 1299 6 1 2 209 1275
0 1300 3 1 2 210 1276
0 1301 6 1 2 146 1277
0 1302 3 1 2 147 1278
0 1303 6 1 2 139 1279
0 1304 3 1 2 140 1280
0 1305 6 1 2 132 1281
0 1306 3 1 2 133 1282
0 1307 6 1 2 125 1283
0 1308 3 1 2 126 1284
0 1309 6 1 2 90 1285
0 1310 3 1 2 91 1286
0 1311 6 1 2 83 1287
0 1312 3 1 2 84 1288
0 1313 6 1 2 76 1289
0 1314 3 1 2 77 1290
0 1315 6 1 2 69 1291
0 1316 3 1 2 70 1292
2 1317 1 1257 
2 1318 1 1257 
2 1319 1 1258 
2 1320 1 1258 
2 1321 1 1259 
2 1322 1 1259 
2 1323 1 1260 
2 1324 1 1260 
3 1325 6 0 2 1294 1293
3 1326 6 0 2 1296 1295
3 1327 6 0 2 1298 1297
3 1328 6 0 2 1300 1299
0 1329 6 1 2 174 1317
0 1330 3 1 2 175 1318
0 1331 6 1 2 167 1319
0 1332 3 1 2 168 1320
0 1333 6 1 2 160 1321
0 1334 3 1 2 161 1322
0 1335 6 1 2 153 1323
0 1336 3 1 2 154 1324
3 1337 6 0 2 1302 1301
3 1338 6 0 2 1304 1303
3 1339 6 0 2 1306 1305
3 1340 6 0 2 1308 1307
3 1341 6 0 2 1310 1309
3 1342 6 0 2 1312 1311
3 1343 6 0 2 1314 1313
3 1344 6 0 2 1316 1315
3 1345 6 0 2 1330 1329
3 1346 6 0 2 1332 1331
3 1347 6 0 2 1334 1333
3 1348 6 0 2 1336 1335
