3	1	0	0	0	
1	5	0	3	0	
1	9	0	2	0	
1	12	0	2	0	
1	15	0	3	0	
1	18	0	72	0	
1	23	0	2	0	
1	26	0	2	0	
1	29	0	2	0	
1	32	0	2	0	
1	35	0	2	0	
1	38	0	20	0	
1	41	0	2	0	
1	44	0	2	0	
1	47	0	2	0	
1	50	0	2	0	
1	53	0	1	0	
1	54	0	1	0	
1	55	0	1	0	
1	56	0	1	0	
1	57	0	1	0	
1	58	0	1	0	
1	59	0	1	0	
1	60	0	1	0	
1	61	0	1	0	
1	62	0	1	0	
1	63	0	1	0	
1	64	0	1	0	
1	65	0	1	0	
1	66	0	2	0	
1	69	0	1	0	
1	70	0	2	0	
1	73	0	1	0	
1	74	0	1	0	
1	75	0	1	0	
1	76	0	1	0	
1	77	0	1	0	
1	78	0	1	0	
1	79	0	1	0	
1	80	0	1	0	
1	81	0	1	0	
1	82	0	1	0	
1	83	0	1	0	
1	84	0	1	0	
1	85	0	1	0	
1	86	0	1	0	
1	87	0	1	0	
1	88	0	1	0	
1	89	0	4	0	
1	94	0	2	0	
1	97	0	2	0	
1	100	0	2	0	
1	103	0	2	0	
3	106	0	0	0	
1	109	0	1	0	
1	110	0	1	0	
1	111	0	1	0	
1	112	0	1	0	
1	113	0	1	0	
1	114	0	1	0	
1	115	0	2	0	
1	118	0	2	0	
1	121	0	2	0	
1	124	0	2	0	
1	127	0	2	0	
1	130	0	2	0	
1	133	0	1	0	
1	134	0	1	0	
1	135	0	2	0	
1	138	0	2	0	
1	141	0	2	0	
1	144	0	2	0	
1	147	0	2	0	
1	150	0	1	0	
1	151	0	1	0	
1	152	0	1	0	
1	153	0	1	0	
1	154	0	1	0	
1	155	0	1	0	
1	156	0	1	0	
1	157	0	1	0	
1	158	0	1	0	
1	159	0	1	0	
1	160	0	1	0	
1	161	0	1	0	
1	162	0	1	0	
1	163	0	1	0	
1	164	0	1	0	
1	165	0	1	0	
1	166	0	1	0	
1	167	0	1	0	
1	168	0	1	0	
1	169	0	1	0	
1	170	0	1	0	
1	171	0	1	0	
1	172	0	1	0	
1	173	0	1	0	
1	174	0	1	0	
1	175	0	1	0	
1	176	0	1	0	
1	177	0	1	0	
1	178	0	1	0	
1	179	0	1	0	
1	180	0	1	0	
1	181	0	1	0	
1	182	0	1	0	
1	183	0	1	0	
1	184	0	1	0	
1	185	0	1	0	
1	186	0	1	0	
1	187	0	1	0	
1	188	0	1	0	
1	189	0	1	0	
1	190	0	1	0	
1	191	0	1	0	
1	192	0	1	0	
1	193	0	1	0	
1	194	0	1	0	
1	195	0	1	0	
1	196	0	1	0	
1	197	0	1	0	
1	198	0	1	0	
1	199	0	1	0	
1	200	0	1	0	
1	201	0	1	0	
1	202	0	1	0	
1	203	0	1	0	
1	204	0	1	0	
1	205	0	1	0	
1	206	0	1	0	
1	207	0	1	0	
1	208	0	1	0	
1	209	0	1	0	
1	210	0	1	0	
1	211	0	1	0	
1	212	0	1	0	
1	213	0	1	0	
1	214	0	1	0	
1	215	0	1	0	
1	216	0	1	0	
1	217	0	1	0	
1	218	0	1	0	
1	219	0	1	0	
1	220	0	1	0	
1	221	0	1	0	
1	222	0	1	0	
1	223	0	1	0	
1	224	0	1	0	
1	225	0	1	0	
1	226	0	1	0	
1	227	0	1	0	
1	228	0	1	0	
1	229	0	1	0	
1	230	0	1	0	
1	231	0	1	0	
1	232	0	1	0	
1	233	0	1	0	
1	234	0	1	0	
1	235	0	1	0	
1	236	0	1	0	
1	237	0	1	0	
1	238	0	1	0	
1	239	0	1	0	
1	240	0	1	0	
3	241	0	0	0	
1	242	0	2	0	
1	245	0	2	0	
3	248	0	0	0	
3	251	0	0	0	
3	254	0	0	0	
3	257	0	0	0	
3	260	0	0	0	
3	263	0	0	0	
3	267	0	0	0	
1	271	0	2	0	
3	274	0	0	0	
3	277	0	0	0	
3	280	0	0	0	
3	283	0	0	0	
3	286	0	0	0	
3	289	0	0	0	
3	293	0	0	0	
3	296	0	0	0	
3	299	0	0	0	
3	303	0	0	0	
3	307	0	0	0	
3	310	0	0	0	
3	313	0	0	0	
3	316	0	0	0	
3	319	0	0	0	
3	322	0	0	0	
3	325	0	0	0	
3	328	0	0	0	
3	331	0	0	0	
3	334	0	0	0	
3	337	0	0	0	
3	340	0	0	0	
3	343	0	0	0	
3	346	0	0	0	
3	349	0	0	0	
3	352	0	0	0	
3	355	0	0	0	
3	358	0	0	0	
3	361	0	0	0	
3	364	0	0	0	
1	367	0	18	0	
1	382	0	4	0	
0	467	5	1	1	57	
0	469	7	2	2	134	133	
0	494	7	2	4	162	172	188	199	
0	528	7	2	4	150	184	228	240	
0	575	7	2	4	183	182	185	186	
0	578	7	2	4	210	152	218	230	
3	582	5	0	1	11356	
0	585	5	1	1	11345	
0	593	5	2	1	11346	
0	596	5	2	1	11347	
0	599	5	6	1	11547	
0	604	5	6	1	11551	
0	609	5	6	1	11553	
0	628	6	13	2	11352	11350	
0	632	6	13	2	11353	11351	
0	641	5	1	1	11531	
0	642	5	1	1	248	
0	644	5	8	1	251	
0	651	5	7	1	254	
0	660	5	7	1	257	
0	666	5	7	1	260	
0	672	5	1	1	11535	
0	673	5	1	1	11537	
0	674	5	1	1	11487	
0	688	7	1	2	11590	11536	
0	695	5	14	1	11361	
0	700	6	6	2	11591	11538	
0	705	5	1	1	11539	
0	706	5	1	1	274	
0	708	5	8	1	277	
0	715	5	7	1	280	
0	721	5	7	1	283	
0	727	5	7	1	286	
0	733	5	1	1	11548	
0	734	5	9	1	293	
0	742	5	7	1	296	
0	748	5	1	1	11552	
0	749	5	1	1	11554	
0	758	5	1	1	307	
0	759	5	2	1	310	
0	762	5	7	1	313	
0	768	5	7	1	316	
0	774	5	7	1	319	
0	780	5	7	1	322	
0	786	5	9	1	325	
0	794	5	7	1	328	
0	800	5	7	1	331	
0	806	5	7	1	334	
0	812	5	1	1	337	
0	814	5	8	1	340	
0	821	5	7	1	343	
0	827	5	7	1	346	
0	833	5	7	1	349	
0	839	5	7	1	352	
0	845	5	9	1	355	
0	853	5	7	1	358	
0	859	5	7	1	361	
0	865	5	7	1	364	
3	881	6	0	2	467	585	
3	882	5	0	1	11600	
3	883	5	0	1	11608	
3	884	5	0	1	11606	
3	885	5	0	1	11598	
0	886	7	1	2	11601	11609	
0	887	7	1	2	11607	11599	
0	957	5	8	1	688	
0	1028	7	1	2	11592	641	
0	1029	6	3	2	11593	705	
0	1109	7	1	2	11596	11612	
3	1110	6	0	2	11529	11610	
3	1111	5	0	1	11357	
3	1112	6	0	2	11530	11611	
3	1113	6	0	2	11597	11613	
3	1114	5	0	1	11358	
0	1115	5	1	1	11570	
0	1167	7	4	2	11716	11443	
0	1174	7	1	2	11717	11444	
0	1189	5	6	1	11488	
0	1194	5	24	1	11362	
0	1199	5	12	1	11363	
0	1206	5	24	1	11364	
0	1218	5	3	1	11571	
0	1222	5	3	1	1028	
3	1489	5	0	1	1109	
0	1537	7	6	2	11967	11445	
0	1551	7	3	2	11446	11968	
0	1649	7	1	2	11993	11447	
0	1708	4	2	2	11969	11448	
0	1721	4	2	2	11449	11970	
3	1781	7	0	2	163	1	
0	1782	7	1	2	170	11365	
0	1783	5	5	1	11366	
0	1789	5	3	1	11367	
0	1793	7	1	2	169	11368	
0	1794	7	1	2	168	11369	
0	1795	7	1	2	167	11370	
0	1796	7	1	2	166	11371	
0	1797	7	1	2	165	11372	
0	1798	7	1	2	164	11373	
0	1799	5	5	1	11374	
0	1805	5	5	1	11375	
0	1811	7	1	2	177	11376	
0	1812	7	1	2	176	11377	
0	1813	7	1	2	175	11378	
0	1814	7	1	2	174	11379	
0	1815	7	1	2	173	11380	
0	1816	7	1	2	157	11381	
0	1817	7	1	2	156	11382	
0	1818	7	1	2	155	11383	
0	1819	7	1	2	154	11384	
0	1820	7	1	2	153	11385	
0	1821	5	1	1	11718	
0	1822	5	1	1	11450	
0	1828	5	1	1	11693	
0	1829	5	1	1	11683	
0	1830	5	1	1	11676	
0	1832	5	1	1	11451	
0	1833	5	1	1	11664	
0	1834	5	1	1	11719	
0	1835	5	1	1	11452	
0	1839	5	1	1	11453	
0	1840	5	1	1	11694	
0	1841	5	1	1	11684	
0	1842	5	1	1	11677	
0	1843	5	1	1	11665	
0	1845	5	5	1	11386	
0	1851	5	5	1	11387	
0	1857	7	1	2	181	11388	
0	1858	7	1	2	171	11389	
0	1859	7	1	2	180	11390	
0	1860	7	1	2	179	11391	
0	1861	7	1	2	178	11392	
0	1862	7	1	2	161	11393	
0	1863	7	1	2	151	11394	
0	1864	7	1	2	160	11395	
0	1865	7	1	2	159	11396	
0	1866	7	1	2	158	11397	
0	1867	5	1	1	11626	
0	1868	5	1	1	11620	
0	1869	5	1	1	11775	
0	1870	5	1	1	11614	
0	1871	5	1	1	11749	
0	1872	5	1	1	11742	
0	1873	5	1	1	11735	
0	1874	5	1	1	11761	
0	1875	5	1	1	11725	
0	1876	5	1	1	11627	
0	1877	5	1	1	11621	
0	1878	5	1	1	11776	
0	1879	5	1	1	11762	
0	1880	5	1	1	11615	
0	1881	5	1	1	11750	
0	1882	5	1	1	11743	
0	1883	5	1	1	11736	
0	1884	5	1	1	11726	
0	1913	5	5	1	11702	
0	1926	7	1	2	11465	11703	
0	1927	7	1	2	11463	11704	
0	1928	7	1	2	11437	11705	
0	1929	7	1	2	11435	11706	
0	1930	7	1	2	11433	11707	
0	1931	5	1	1	11858	
0	1932	5	1	1	11849	
0	1933	5	1	1	11842	
0	1934	5	1	1	11827	
0	1935	5	1	1	11820	
0	1936	5	1	1	11811	
0	1937	5	1	1	11804	
0	1938	5	1	1	11795	
0	1939	5	1	1	11859	
0	1940	5	1	1	11850	
0	1941	5	1	1	11843	
0	1942	5	1	1	11821	
0	1943	5	1	1	11812	
0	1944	5	1	1	11805	
0	1945	5	1	1	11796	
0	1946	5	1	1	11828	
0	1947	5	5	1	11398	
0	1953	5	3	1	11399	
0	1957	7	1	2	209	11400	
0	1958	7	1	2	216	11401	
0	1959	7	1	2	215	11402	
0	1960	7	1	2	214	11403	
0	1961	7	1	2	213	11404	
0	1962	7	1	2	212	11405	
0	1963	7	1	2	211	11406	
0	1965	5	1	1	11454	
0	1966	7	1	2	12116	11455	
0	1967	5	1	1	11456	
0	1968	5	1	1	11934	
0	1969	5	1	1	11927	
0	1970	5	1	1	11920	
0	1971	5	1	1	11911	
0	1972	5	1	1	11902	
0	1973	5	1	1	11892	
0	1974	5	1	1	11885	
0	1975	5	1	1	11878	
0	1976	5	1	1	11870	
0	1977	5	5	1	11407	
0	1983	5	5	1	11408	
0	1989	7	1	2	642	11409	
0	1990	7	1	2	11666	11410	
0	1991	7	1	2	11678	11411	
0	1992	7	1	2	674	11412	
0	1993	7	1	2	11685	11413	
0	1994	7	1	2	11695	11414	
0	1995	7	1	2	672	11415	
0	1996	7	1	2	673	11416	
0	1997	5	5	1	11708	
0	2010	7	1	2	11467	11709	
0	2011	7	1	2	11441	11710	
0	2012	7	1	2	11439	11711	
0	2013	7	1	2	11469	11712	
0	2014	7	1	2	11471	11713	
0	2015	5	1	1	11935	
0	2016	5	1	1	11928	
0	2017	5	1	1	11921	
0	2018	5	1	1	11903	
0	2019	5	1	1	11893	
0	2020	5	1	1	11886	
0	2021	5	1	1	11879	
0	2022	5	1	1	11912	
0	2023	5	1	1	11871	
0	2052	5	5	1	11417	
0	2058	5	5	1	11418	
0	2064	7	1	2	706	11419	
0	2065	7	1	2	11727	11420	
0	2066	7	1	2	11737	11421	
0	2067	7	1	2	11744	11422	
0	2068	7	1	2	11751	11423	
0	2069	7	1	2	733	11424	
0	2070	7	1	2	11763	11425	
0	2071	7	1	2	11777	11426	
0	2072	7	1	2	748	11427	
0	2073	7	1	2	749	11428	
0	2107	6	1	2	11457	1821	
0	2108	6	1	2	11720	1822	
0	2110	5	1	1	11971	
0	2111	6	1	2	11972	1832	
0	2112	6	1	2	11458	1834	
0	2113	6	1	2	11721	1835	
0	2114	5	1	1	11973	
0	2115	6	1	2	11974	1839	
0	2117	5	1	1	12251	
0	2171	5	1	1	11994	
0	2172	6	1	2	11995	1965	
0	2230	5	1	1	12249	
0	2239	3	1	2	12273	1782	
0	2240	3	1	2	12274	11429	
0	2241	3	1	2	12275	1793	
0	2242	3	1	2	12276	1794	
0	2243	3	1	2	12277	1795	
0	2244	3	1	2	12278	1796	
0	2245	3	1	2	12279	1797	
0	2246	3	1	2	12280	1798	
0	2247	3	1	2	12283	1811	
0	2248	3	1	2	12284	1812	
0	2249	3	1	2	12285	1813	
0	2250	3	1	2	12286	1814	
0	2251	3	1	2	12287	1815	
0	2252	3	1	2	12296	1816	
0	2253	3	1	2	12297	1817	
0	2254	3	1	2	12298	1818	
0	2255	3	1	2	12299	1819	
0	2256	3	1	2	12300	1820	
0	2257	6	11	2	2107	2108	
0	2267	5	1	1	12038	
0	2268	6	1	2	11459	2110	
0	2269	6	6	2	2112	2113	
0	2274	6	1	2	11460	2114	
0	2275	5	1	1	12039	
0	2277	7	1	2	11518	12307	
0	2278	7	1	2	11525	12308	
0	2279	7	1	2	11509	12309	
0	2280	7	1	2	11523	12310	
0	2281	7	1	2	11507	12311	
0	2282	7	1	2	11519	12312	
0	2283	7	1	2	11526	12313	
0	2284	7	1	2	11510	12314	
0	2285	7	1	2	11524	12315	
0	2286	7	1	2	11508	12316	
0	2287	5	5	1	12074	
0	2293	5	5	1	12044	
0	2299	7	1	2	11485	12075	
0	2300	7	1	2	11505	12076	
0	2301	7	1	2	11503	12077	
0	2302	7	1	2	11501	12078	
0	2303	7	1	2	11483	12079	
0	2304	7	1	2	11486	12045	
0	2305	7	1	2	11506	12046	
0	2306	7	1	2	11504	12047	
0	2307	7	1	2	11502	12048	
0	2308	7	1	2	11484	12049	
0	2309	5	5	1	12080	
0	2315	5	5	1	12050	
0	2321	7	1	2	11489	12081	
0	2322	7	1	2	11497	12082	
0	2323	7	1	2	11481	12083	
0	2324	7	1	2	11479	12084	
0	2325	7	1	2	11499	12085	
0	2326	7	1	2	11490	12051	
0	2327	7	1	2	11498	12052	
0	2328	7	1	2	11482	12053	
0	2329	7	1	2	11480	12054	
0	2330	7	1	2	11500	12055	
0	2331	5	5	1	12056	
0	2337	7	1	2	208	12321	
0	2338	7	1	2	198	12322	
0	2339	7	1	2	207	12323	
0	2340	7	1	2	206	12324	
0	2341	7	1	2	205	12325	
0	2342	7	1	2	11466	12057	
0	2343	7	1	2	11464	12058	
0	2344	7	1	2	11438	12059	
0	2345	7	1	2	11436	12060	
0	2346	7	1	2	11434	12061	
0	2347	3	1	2	12331	11430	
0	2348	3	1	2	12332	1957	
0	2349	3	1	2	12333	1958	
0	2350	3	1	2	12334	1959	
0	2351	3	1	2	12335	1960	
0	2352	3	1	2	12336	1961	
0	2353	3	1	2	12337	1962	
0	2354	3	1	2	12338	1963	
0	2355	6	1	2	11461	2171	
0	2356	5	1	1	12117	
0	2357	6	1	2	12118	1967	
0	2358	7	1	2	114	12346	
0	2359	7	1	2	113	12347	
0	2360	7	1	2	111	12348	
0	2361	7	1	2	87	12349	
0	2362	7	1	2	112	12350	
0	2363	7	1	2	88	12351	
0	2364	7	1	2	11532	12352	
0	2365	7	1	2	11540	12353	
0	2366	7	1	2	11790	12354	
0	2367	7	1	2	11473	12355	
0	2368	5	5	1	12062	
0	2374	7	1	2	193	12360	
0	2375	7	1	2	192	12361	
0	2376	7	1	2	191	12362	
0	2377	7	1	2	190	12363	
0	2378	7	1	2	189	12364	
0	2379	7	1	2	11468	12063	
0	2380	7	1	2	11442	12064	
0	2381	7	1	2	11440	12065	
0	2382	7	1	2	11470	12066	
0	2383	7	1	2	11472	12067	
0	2384	5	5	1	12086	
0	2390	5	5	1	12087	
0	2396	7	1	2	58	12088	
0	2397	7	1	2	77	12089	
0	2398	7	1	2	78	12090	
0	2399	7	1	2	59	12091	
0	2400	7	1	2	81	12092	
0	2401	7	1	2	80	12093	
0	2402	7	1	2	79	12094	
0	2403	7	1	2	60	12095	
0	2404	7	1	2	61	12096	
0	2405	7	1	2	62	12097	
0	2406	5	5	1	12098	
0	2412	5	5	1	12099	
0	2418	7	1	2	69	12100	
0	2419	7	1	2	11474	12101	
0	2420	7	1	2	74	12102	
0	2421	7	1	2	76	12103	
0	2422	7	1	2	75	12104	
0	2423	7	1	2	73	12105	
0	2424	7	1	2	53	12106	
0	2425	7	1	2	54	12107	
0	2426	7	1	2	55	12108	
0	2427	7	1	2	56	12109	
0	2428	7	1	2	82	12377	
0	2429	7	1	2	65	12378	
0	2430	7	1	2	83	12379	
0	2431	7	1	2	84	12380	
0	2432	7	1	2	85	12381	
0	2433	7	1	2	64	12382	
0	2434	7	1	2	63	12383	
0	2435	7	1	2	86	12384	
0	2436	7	1	2	109	12385	
0	2437	7	1	2	110	12386	
0	2441	7	1	2	2239	11638	
0	2442	7	5	2	2240	11639	
0	2446	7	5	2	2241	11640	
0	2450	7	5	2	2242	11641	
0	2454	7	5	2	2243	11642	
0	2458	7	5	2	2244	11643	
0	2462	7	5	2	2247	11644	
0	2466	7	5	2	2248	11645	
0	2470	7	5	2	2249	11646	
0	2474	7	5	2	2250	11647	
0	2478	7	5	2	2251	11648	
0	2482	7	8	2	2252	11651	
0	2488	7	10	2	2253	11652	
0	2496	7	8	2	2254	11653	
0	2502	7	8	2	2255	11654	
0	2508	7	8	2	2256	11655	
0	2523	6	7	2	2268	2111	
0	2533	6	3	2	2274	2115	
0	2537	5	1	1	12218	
0	2538	3	5	2	2278	1858	
0	2542	3	5	2	2279	1859	
0	2546	3	5	2	2280	1860	
0	2550	3	5	2	2281	1861	
0	2554	3	9	2	2283	1863	
0	2561	3	8	2	2284	1864	
0	2567	3	8	2	2285	1865	
0	2573	3	8	2	2286	1866	
0	2604	3	3	2	2338	1927	
0	2607	3	5	2	2339	1928	
0	2611	3	5	2	2340	1929	
0	2615	3	5	2	2341	1930	
0	2619	7	9	2	2348	11656	
0	2626	7	8	2	2349	11657	
0	2632	7	8	2	2350	11658	
0	2638	7	8	2	2351	11659	
0	2644	7	8	2	2352	11660	
0	2650	6	2	2	2355	2172	
0	2653	6	1	2	11462	2356	
0	2654	3	5	2	2359	1990	
0	2658	3	5	2	2360	1991	
0	2662	3	5	2	2361	1992	
0	2666	3	5	2	2362	1993	
0	2670	3	5	2	2363	1994	
0	2674	3	7	2	2366	11431	
0	2680	3	3	2	2367	11432	
0	2688	3	5	2	2374	2010	
0	2692	3	5	2	2375	2011	
0	2696	3	5	2	2376	2012	
0	2700	3	5	2	2377	2013	
0	2704	3	5	2	2378	2014	
0	2728	7	1	2	2347	11661	
0	2729	3	5	2	2429	2065	
0	2733	3	5	2	2430	2066	
0	2737	3	5	2	2431	2067	
0	2741	3	5	2	2432	2068	
0	2745	3	5	2	2433	2069	
0	2749	3	5	2	2434	2070	
0	2753	3	5	2	2435	2071	
0	2757	3	5	2	2436	2072	
0	2761	3	5	2	2437	2073	
0	2765	5	1	1	12212	
0	2766	7	2	2	2354	11662	
0	2769	7	2	2	2353	11663	
0	2772	7	2	2	2246	11649	
0	2775	7	2	2	2245	11650	
0	2778	3	2	2	2282	1862	
0	2781	3	2	2	2358	1989	
0	2784	3	2	2	2365	1996	
0	2787	3	2	2	2364	1995	
0	2790	3	2	2	2337	1926	
0	2793	3	2	2	2277	1857	
0	2796	3	2	2	2428	2064	
0	2866	7	1	2	12454	12213	
0	2867	7	1	2	12455	12214	
0	2868	7	1	2	12456	12215	
0	2869	7	1	2	12457	12216	
0	2878	7	1	2	12465	12219	
0	2913	7	1	2	204	12471	
0	2914	7	1	2	203	12472	
0	2915	7	1	2	202	12473	
0	2916	7	1	2	201	12474	
0	2917	7	1	2	200	12475	
0	2918	7	1	2	235	12479	
0	2919	7	1	2	234	12480	
0	2920	7	1	2	233	12481	
0	2921	7	1	2	232	12482	
0	2922	7	1	2	231	12483	
0	2923	7	1	2	197	12484	
0	2924	7	1	2	187	12485	
0	2925	7	1	2	196	12486	
0	2926	7	1	2	195	12487	
0	2927	7	1	2	194	12488	
0	2928	7	1	2	227	12492	
0	2929	7	1	2	217	12493	
0	2930	7	1	2	226	12494	
0	2931	7	1	2	225	12495	
0	2932	7	1	2	224	12496	
0	2933	7	1	2	239	12501	
0	2934	7	1	2	229	12502	
0	2935	7	1	2	238	12503	
0	2936	7	1	2	237	12504	
0	2937	7	1	2	236	12505	
0	2988	6	1	2	2653	2357	
0	3005	7	1	2	223	12508	
0	3006	7	1	2	222	12509	
0	3007	7	1	2	221	12510	
0	3008	7	1	2	220	12511	
0	3009	7	1	2	219	12512	
0	3020	7	1	2	812	12513	
0	3021	7	1	2	11872	12514	
0	3022	7	1	2	11880	12515	
0	3023	7	1	2	11887	12516	
0	3024	7	1	2	11894	12517	
0	3025	7	1	2	11904	12518	
0	3026	7	1	2	11913	12519	
0	3027	7	1	2	11922	12520	
0	3028	7	1	2	11929	12521	
0	3029	7	1	2	11936	12522	
0	3032	7	1	2	758	12523	
0	3033	7	1	2	11791	12524	
0	3034	7	1	2	11797	12525	
0	3035	7	1	2	11806	12526	
0	3036	7	1	2	11813	12527	
0	3037	7	1	2	11822	12528	
0	3038	7	1	2	11829	12529	
0	3039	7	1	2	11844	12530	
0	3040	7	1	2	11851	12531	
0	3041	7	1	2	11860	12532	
0	3073	5	2	1	2728	
0	3080	5	2	1	2441	
0	3096	7	1	2	11696	12786	
0	3097	7	3	2	11686	12778	
0	3101	7	5	2	12040	12770	
0	3107	7	6	2	11679	12760	
0	3114	7	8	2	11667	12747	
0	3122	7	3	2	12648	12458	
0	3126	3	3	2	12034	2866	
0	3130	7	1	2	12649	12459	
0	3131	3	2	2	12035	2869	
0	3134	7	1	2	12650	12460	
0	3135	5	1	1	12655	
0	3136	7	1	2	11697	12787	
0	3137	7	2	2	11687	12779	
0	3140	7	3	2	12041	12771	
0	3144	7	4	2	11680	12761	
0	3149	7	5	2	11668	12748	
0	3155	7	3	2	12656	12466	
0	3159	3	3	2	1174	2878	
0	3167	5	1	1	12937	
0	3168	7	1	2	11628	12638	
0	3169	7	3	2	11622	12628	
0	3173	7	4	2	11778	12618	
0	3178	7	6	2	11764	12608	
0	3184	7	1	2	11616	12596	
0	3185	7	3	2	11752	12705	
0	3189	7	5	2	11745	12697	
0	3195	7	6	2	11738	12689	
0	3202	7	8	2	11728	12680	
0	3210	7	1	2	11629	12639	
0	3211	7	3	2	11623	12629	
0	3215	7	5	2	11779	12619	
0	3221	7	7	2	12609	11765	
0	3228	7	1	2	11617	12597	
0	3229	7	2	2	11753	12706	
0	3232	7	3	2	11746	12698	
0	3236	7	4	2	11739	12690	
0	3241	7	5	2	11729	12681	
0	3247	3	5	2	2913	2299	
0	3251	3	5	2	2914	2300	
0	3255	3	5	2	2915	2301	
0	3259	3	5	2	2916	2302	
0	3263	3	5	2	2917	2303	
0	3267	3	8	2	2918	2304	
0	3273	3	10	2	2919	2305	
0	3281	3	8	2	2920	2306	
0	3287	3	8	2	2921	2307	
0	3293	3	8	2	2922	2308	
0	3299	3	5	2	2924	2322	
0	3303	3	5	2	2925	2323	
0	3307	3	5	2	2926	2324	
0	3311	3	5	2	2927	2325	
0	3315	3	9	2	2929	2327	
0	3322	3	8	2	2930	2328	
0	3328	3	8	2	2931	2329	
0	3334	3	8	2	2932	2330	
0	3340	3	3	2	2934	2343	
0	3343	3	8	2	2935	2344	
0	3349	3	8	2	2936	2345	
0	3355	3	8	2	2937	2346	
0	3361	7	1	2	12920	12591	
0	3362	7	1	2	12913	12584	
0	3363	7	1	2	12906	12575	
0	3364	7	1	2	12897	12568	
0	3365	7	1	2	12890	12558	
0	3366	7	1	2	12885	12675	
0	3367	7	1	2	12878	12668	
0	3368	7	1	2	12871	12663	
0	3369	7	1	2	12866	12658	
0	3370	7	1	2	12816	12553	
0	3371	7	1	2	12811	12548	
0	3372	7	1	2	12806	12543	
0	3373	7	1	2	12801	12538	
0	3374	7	1	2	12796	12533	
0	3375	7	3	2	2988	12794	
0	3379	7	1	2	12795	1966	
0	3380	5	1	1	12939	
0	3381	7	3	2	11714	12721	
0	3384	3	8	2	3005	2379	
0	3390	3	10	2	3006	2380	
0	3398	3	8	2	3007	2381	
0	3404	3	8	2	3008	2382	
0	3410	3	8	2	3009	2383	
0	3416	3	5	2	3021	2397	
0	3420	3	5	2	3022	2398	
0	3424	3	5	2	3023	2399	
0	3428	3	5	2	3024	2400	
0	3432	3	5	2	3025	2401	
0	3436	3	5	2	3026	2402	
0	3440	3	5	2	3027	2403	
0	3444	3	5	2	3028	2404	
0	3448	3	5	2	3029	2405	
0	3452	5	1	1	12945	
0	3453	5	1	1	12947	
0	3454	3	5	2	3034	2420	
0	3458	3	5	2	3035	2421	
0	3462	3	5	2	3036	2422	
0	3466	3	5	2	3037	2423	
0	3470	3	5	2	3038	2424	
0	3474	3	5	2	3039	2425	
0	3478	3	5	2	3040	2426	
0	3482	3	5	2	3041	2427	
0	3486	5	1	1	12949	
0	3507	4	2	2	12036	2868	
0	3515	4	2	2	11669	12749	
0	3551	5	1	1	12927	
0	3552	5	1	1	12931	
0	3569	5	1	1	12933	
0	3570	5	1	1	12935	
0	3625	4	2	2	11766	12610	
0	3628	4	2	2	11730	12682	
0	3658	4	2	2	12611	11767	
0	3781	5	1	1	12941	
0	3782	5	1	1	12943	
0	3783	3	2	2	2928	2326	
0	3786	3	2	2	2933	2342	
0	3789	3	2	2	2923	2321	
0	3885	3	2	2	3033	2419	
0	3888	3	2	2	3032	2418	
0	3891	3	2	2	3020	2396	
0	3953	6	1	2	12467	2117	
0	3954	5	1	1	12468	
0	3955	6	1	2	12469	2537	
0	3956	5	1	1	12470	
0	3958	5	1	1	13019	
0	3964	5	1	1	13021	
0	4193	3	3	2	1649	3379	
0	4303	3	2	3	12037	2867	3130	
0	4308	5	1	1	12461	
0	4313	5	1	1	12462	
0	4326	6	1	2	12932	3551	
0	4327	6	1	2	12928	3552	
0	4333	6	1	2	12936	3569	
0	4334	6	1	2	12934	3570	
0	4411	6	1	2	12944	3781	
0	4412	6	1	2	12942	3782	
0	4463	6	1	2	12788	1828	
0	4464	5	1	1	12789	
0	4465	6	1	2	12780	1829	
0	4466	5	1	1	12781	
0	4467	6	1	2	12772	2267	
0	4468	5	1	1	12773	
0	4469	6	1	2	12762	1830	
0	4470	5	1	1	12763	
0	4471	6	1	2	12750	1833	
0	4472	5	1	1	12751	
0	4473	5	1	1	13051	
0	4474	5	1	1	13054	
0	4475	6	1	2	12790	1840	
0	4476	5	1	1	12791	
0	4477	6	1	2	12782	1841	
0	4478	5	1	1	12783	
0	4479	6	1	2	12774	2275	
0	4480	5	1	1	12775	
0	4481	6	1	2	12764	1842	
0	4482	5	1	1	12765	
0	4483	6	1	2	12752	1843	
0	4484	5	1	1	12753	
0	4485	5	1	1	13077	
0	4486	5	1	1	13080	
0	4487	6	1	2	12252	3954	
0	4488	6	1	2	12220	3956	
0	4489	5	1	1	12754	
0	4490	6	1	2	12755	3958	
0	4491	5	1	1	12776	
0	4492	5	1	1	12766	
0	4493	5	1	1	12792	
0	4494	5	1	1	12784	
0	4495	5	1	1	12534	
0	4496	6	1	2	12535	3964	
0	4497	5	1	1	12544	
0	4498	5	1	1	12539	
0	4499	5	1	1	12554	
0	4500	5	1	1	12549	
0	4501	5	1	1	12683	
0	4502	6	1	2	12684	3167	
0	4503	5	1	1	12699	
0	4504	5	1	1	12691	
0	4505	5	1	1	12598	
0	4506	5	1	1	12707	
0	4507	6	1	2	12640	1867	
0	4508	5	1	1	12641	
0	4509	6	1	2	12630	1868	
0	4510	5	1	1	12631	
0	4511	6	1	2	12620	1869	
0	4512	5	1	1	12621	
0	4513	6	1	2	12599	1870	
0	4514	5	1	1	12600	
0	4515	6	1	2	12708	1871	
0	4516	5	1	1	12709	
0	4517	6	1	2	12700	1872	
0	4518	5	1	1	12701	
0	4519	6	1	2	12692	1873	
0	4520	5	1	1	12693	
0	4521	6	1	2	12612	1874	
0	4522	5	1	1	12613	
0	4523	6	1	2	12685	1875	
0	4524	5	1	1	12686	
0	4525	6	1	2	12642	1876	
0	4526	5	1	1	12643	
0	4527	6	1	2	12632	1877	
0	4528	5	1	1	12633	
0	4529	6	1	2	12622	1878	
0	4530	5	1	1	12623	
0	4531	6	1	2	12614	1879	
0	4532	5	1	1	12615	
0	4533	6	1	2	12601	1880	
0	4534	5	1	1	12602	
0	4535	6	1	2	12710	1881	
0	4536	5	1	1	12711	
0	4537	6	1	2	12702	1882	
0	4538	5	1	1	12703	
0	4539	6	1	2	12694	1883	
0	4540	5	1	1	12695	
0	4541	6	1	2	12687	1884	
0	4542	5	1	1	12688	
0	4543	5	1	1	13435	
0	4544	7	1	2	11861	13206	
0	4545	7	3	2	11852	13198	
0	4549	7	5	2	11845	13190	
0	4555	7	7	2	13180	11830	
0	4562	7	1	2	11823	13172	
0	4563	7	2	2	11814	13286	
0	4566	7	3	2	11807	13278	
0	4570	7	4	2	11798	13270	
0	4575	5	1	1	12821	
0	4576	7	1	2	11862	13207	
0	4577	7	3	2	11853	13199	
0	4581	7	4	2	11846	13191	
0	4586	7	6	2	11831	13181	
0	4592	7	1	2	11824	13173	
0	4593	7	3	2	11815	13287	
0	4597	7	5	2	11808	13279	
0	4603	7	6	2	11799	13271	
0	4610	5	1	1	12822	
0	4611	5	1	1	12921	
0	4612	5	1	1	12592	
0	4613	5	1	1	12914	
0	4614	5	1	1	12585	
0	4615	5	1	1	12907	
0	4616	5	1	1	12576	
0	4617	5	1	1	12891	
0	4618	5	1	1	12559	
0	4619	5	1	1	12886	
0	4620	5	1	1	12676	
0	4621	5	1	1	12879	
0	4622	5	1	1	12669	
0	4623	5	1	1	12872	
0	4624	5	1	1	12664	
0	4625	5	1	1	12898	
0	4626	5	1	1	12569	
0	4627	5	1	1	12867	
0	4628	5	1	1	12659	
0	4629	5	1	1	12857	
0	4630	7	1	2	13382	12858	
0	4631	5	1	1	12850	
0	4632	7	1	2	13377	12851	
0	4633	5	1	1	12845	
0	4634	7	1	2	13372	12846	
0	4635	7	1	2	13367	12840	
0	4636	5	1	1	12833	
0	4637	7	1	2	13362	12834	
0	4638	7	1	2	13357	13229	
0	4639	7	1	2	13352	13224	
0	4640	7	1	2	13347	13219	
0	4641	7	1	2	13342	13214	
0	4642	5	1	1	12841	
0	4643	5	1	1	12817	
0	4644	5	1	1	12555	
0	4645	5	1	1	12812	
0	4646	5	1	1	12550	
0	4647	5	1	1	12807	
0	4648	5	1	1	12545	
0	4649	5	1	1	12802	
0	4650	5	1	1	12540	
0	4651	5	1	1	12797	
0	4652	5	1	1	12536	
0	4653	5	1	1	13294	
0	4656	7	1	2	11937	13334	
0	4657	7	3	2	11930	13326	
0	4661	7	5	2	11923	13318	
0	4667	7	7	2	13308	11914	
0	4674	7	1	2	11905	13300	
0	4675	7	2	2	11895	13259	
0	4678	7	3	2	11888	13251	
0	4682	7	4	2	11881	13243	
0	4687	7	5	2	11873	13234	
0	4693	5	1	1	12798	
0	4694	6	1	2	12799	3380	
0	4695	5	1	1	12808	
0	4696	5	1	1	12803	
0	4697	5	1	1	12818	
0	4698	5	1	1	12813	
0	4699	5	1	1	13437	
0	4700	5	1	1	13439	
0	4701	7	1	2	11938	13335	
0	4702	7	3	2	11931	13327	
0	4706	7	4	2	11924	13319	
0	4711	7	6	2	11915	13309	
0	4717	7	1	2	11906	13301	
0	4718	7	3	2	11896	13260	
0	4722	7	5	2	11889	13252	
0	4728	7	6	2	11882	13244	
0	4735	7	8	2	11874	13235	
0	4743	5	1	1	13443	
0	4744	5	1	1	12835	
0	4745	5	1	1	12722	
0	4746	6	1	2	12723	3452	
0	4747	5	1	1	12731	
0	4748	5	1	1	12724	
0	4749	5	1	1	12740	
0	4750	5	1	1	12660	
0	4751	6	1	2	12661	3453	
0	4752	5	1	1	12670	
0	4753	5	1	1	12665	
0	4754	5	1	1	12560	
0	4755	5	1	1	12677	
0	4756	7	1	2	13422	13167	
0	4757	7	1	2	13417	13162	
0	4758	7	1	2	13412	13157	
0	4759	7	1	2	13407	13152	
0	4760	7	1	2	13402	13147	
0	4761	5	1	1	12741	
0	4762	7	1	2	13397	12742	
0	4763	5	1	1	12732	
0	4764	7	1	2	13392	12733	
0	4765	5	1	1	12725	
0	4766	7	1	2	13387	12726	
0	4767	7	1	2	12828	13297	
0	4768	5	1	1	12829	
0	4769	7	7	2	13267	11715	
0	4775	5	1	1	12868	
0	4776	6	1	2	12869	3486	
0	4777	5	1	1	12880	
0	4778	5	1	1	12873	
0	4779	5	1	1	12892	
0	4780	5	1	1	12887	
0	4781	5	1	1	13455	
0	4782	5	1	1	13457	
0	4783	5	1	1	13459	
0	4784	3	2	2	13059	3134	
0	4789	5	1	1	12651	
0	4790	5	2	1	13060	
0	4793	5	1	1	13427	
0	4794	5	1	1	12652	
0	4795	5	1	1	13429	
0	4799	5	1	1	12624	
0	4800	5	1	1	12616	
0	4801	5	1	1	12644	
0	4802	5	1	1	12634	
0	4803	6	2	2	4326	4327	
0	4806	6	2	2	4333	4334	
0	4809	5	1	1	13431	
0	4813	5	1	1	13433	
0	4844	4	2	2	13182	11832	
0	4871	4	2	2	11833	13183	
0	4940	4	2	2	13310	11916	
0	4997	6	2	2	4411	4412	
0	5027	4	2	2	11917	13311	
0	5030	4	2	2	11875	13236	
0	5045	5	1	1	12847	
0	5046	5	1	1	12842	
0	5047	5	1	1	12859	
0	5048	5	1	1	12852	
0	5064	5	1	1	12577	
0	5065	5	1	1	12570	
0	5066	5	1	1	12593	
0	5067	5	1	1	12586	
0	5110	5	1	1	12908	
0	5111	5	1	1	12899	
0	5112	5	1	1	12922	
0	5113	5	1	1	12915	
0	5165	6	1	2	4486	4485	
0	5166	6	1	2	4474	4473	
0	5167	6	1	2	11698	4464	
0	5168	6	1	2	11688	4466	
0	5169	6	1	2	12042	4468	
0	5170	6	1	2	11681	4470	
0	5171	6	1	2	11670	4472	
0	5172	6	1	2	11699	4476	
0	5173	6	1	2	11689	4478	
0	5174	6	1	2	12043	4480	
0	5175	6	1	2	11682	4482	
0	5176	6	1	2	11671	4484	
0	5177	6	1	2	3953	4487	
0	5178	6	1	2	3955	4488	
0	5179	6	1	2	13020	4489	
0	5180	6	1	2	12767	4491	
0	5181	6	1	2	12777	4492	
0	5182	6	1	2	12785	4493	
0	5183	6	1	2	12793	4494	
0	5184	6	1	2	13022	4495	
0	5185	6	1	2	12541	4497	
0	5186	6	1	2	12546	4498	
0	5187	6	1	2	12551	4499	
0	5188	6	1	2	12556	4500	
0	5189	6	1	2	12938	4501	
0	5190	6	1	2	12696	4503	
0	5191	6	1	2	12704	4504	
0	5192	6	1	2	12712	4505	
0	5193	6	1	2	12603	4506	
0	5196	6	1	2	11630	4508	
0	5197	6	1	2	11624	4510	
0	5198	6	1	2	11780	4512	
0	5199	6	1	2	11618	4514	
0	5200	6	1	2	11754	4516	
0	5201	6	1	2	11747	4518	
0	5202	6	1	2	11740	4520	
0	5203	6	1	2	11768	4522	
0	5204	6	1	2	11731	4524	
0	5205	6	1	2	11631	4526	
0	5206	6	1	2	11625	4528	
0	5207	6	1	2	11781	4530	
0	5208	6	1	2	11769	4532	
0	5209	6	1	2	11619	4534	
0	5210	6	1	2	11755	4536	
0	5211	6	1	2	11748	4538	
0	5212	6	1	2	11741	4540	
0	5213	6	1	2	11732	4542	
0	5283	6	1	2	12594	4611	
0	5284	6	1	2	12923	4612	
0	5285	6	1	2	12587	4613	
0	5286	6	1	2	12916	4614	
0	5287	6	1	2	12578	4615	
0	5288	6	1	2	12909	4616	
0	5289	6	1	2	12561	4617	
0	5290	6	1	2	12893	4618	
0	5291	6	1	2	12678	4619	
0	5292	6	1	2	12888	4620	
0	5293	6	1	2	12671	4621	
0	5294	6	1	2	12881	4622	
0	5295	6	1	2	12666	4623	
0	5296	6	1	2	12874	4624	
0	5297	6	1	2	12571	4625	
0	5298	6	1	2	12900	4626	
0	5299	6	1	2	12662	4627	
0	5300	6	1	2	12870	4628	
0	5314	6	1	2	12557	4643	
0	5315	6	1	2	12819	4644	
0	5316	6	1	2	12552	4645	
0	5317	6	1	2	12814	4646	
0	5318	6	1	2	12547	4647	
0	5319	6	1	2	12809	4648	
0	5320	6	1	2	12542	4649	
0	5321	6	1	2	12804	4650	
0	5322	6	1	2	12537	4651	
0	5323	6	1	2	12800	4652	
0	5324	5	1	1	13468	
0	5363	6	1	2	12940	4693	
0	5364	6	1	2	12805	4695	
0	5365	6	1	2	12810	4696	
0	5366	6	1	2	12815	4697	
0	5367	6	1	2	12820	4698	
0	5425	6	1	2	12946	4745	
0	5426	6	1	2	12727	4747	
0	5427	6	1	2	12734	4748	
0	5429	6	1	2	12948	4750	
0	5430	6	1	2	12667	4752	
0	5431	6	1	2	12672	4753	
0	5432	6	1	2	12679	4754	
0	5433	6	1	2	12562	4755	
0	5451	6	1	2	12950	4775	
0	5452	6	1	2	12875	4777	
0	5453	6	1	2	12882	4778	
0	5454	6	1	2	12889	4779	
0	5455	6	1	2	12894	4780	
0	5456	6	1	2	13458	4781	
0	5457	6	1	2	13456	4782	
0	5469	5	1	1	13471	
0	5474	6	1	2	12617	4799	
0	5475	6	1	2	12625	4800	
0	5476	6	1	2	12635	4801	
0	5477	6	1	2	12645	4802	
0	5571	6	1	2	12843	5045	
0	5572	6	1	2	12848	5046	
0	5573	6	1	2	12853	5047	
0	5574	6	1	2	12860	5048	
0	5584	6	1	2	12572	5064	
0	5585	6	1	2	12579	5065	
0	5586	6	1	2	12588	5066	
0	5587	6	1	2	12595	5067	
0	5602	6	1	2	12901	5110	
0	5603	6	1	2	12910	5111	
0	5604	6	1	2	12917	5112	
0	5605	6	1	2	12924	5113	
0	5631	6	1	2	5324	4653	
0	5632	6	9	2	4463	5167	
0	5640	6	15	2	4465	5168	
0	5654	6	17	2	4467	5169	
0	5670	6	14	2	4469	5170	
0	5683	6	8	2	4471	5171	
0	5690	6	7	2	4475	5172	
0	5697	6	10	2	4477	5173	
0	5707	6	11	2	4479	5174	
0	5718	6	10	2	4481	5175	
0	5728	6	7	2	4483	5176	
0	5735	5	1	1	5177	
0	5736	6	3	2	5179	4490	
0	5740	6	3	2	5180	5181	
0	5744	6	4	2	5182	5183	
0	5747	6	3	2	5184	4496	
0	5751	6	3	2	5185	5186	
0	5755	6	4	2	5187	5188	
0	5758	6	3	2	5189	4502	
0	5762	6	3	2	5190	5191	
0	5766	6	4	2	5192	5193	
0	5769	5	1	1	13599	
0	5770	5	1	1	13601	
0	5771	6	8	2	4507	5196	
0	5778	6	12	2	4509	5197	
0	5789	6	11	2	4511	5198	
0	5799	6	9	2	4513	5199	
0	5807	6	15	2	4515	5200	
0	5821	6	17	2	4517	5201	
0	5837	6	14	2	4519	5202	
0	5850	6	7	2	4521	5203	
0	5856	6	8	2	4523	5204	
0	5863	6	8	2	4525	5205	
0	5870	6	12	2	4527	5206	
0	5881	6	12	2	4529	5207	
0	5892	6	5	2	4531	5208	
0	5898	6	7	2	4533	5209	
0	5905	6	10	2	4535	5210	
0	5915	6	11	2	4537	5211	
0	5926	6	10	2	4539	5212	
0	5936	6	7	2	4541	5213	
0	5943	5	1	1	13126	
0	5944	6	1	2	13208	1931	
0	5945	5	1	1	13209	
0	5946	6	1	2	13200	1932	
0	5947	5	1	1	13201	
0	5948	6	1	2	13192	1933	
0	5949	5	1	1	13193	
0	5950	6	1	2	13184	1934	
0	5951	5	1	1	13185	
0	5952	6	1	2	13174	1935	
0	5953	5	1	1	13175	
0	5954	6	1	2	13288	1936	
0	5955	5	1	1	13289	
0	5956	6	1	2	13280	1937	
0	5957	5	1	1	13281	
0	5958	6	1	2	13272	1938	
0	5959	5	1	1	13273	
0	5960	7	5	2	12823	13588	
0	5966	5	1	1	13603	
0	5967	6	1	2	13210	1939	
0	5968	5	1	1	13211	
0	5969	6	1	2	13202	1940	
0	5970	5	1	1	13203	
0	5971	6	1	2	13194	1941	
0	5972	5	1	1	13195	
0	5973	6	1	2	13176	1942	
0	5974	5	1	1	13177	
0	5975	6	1	2	13290	1943	
0	5976	5	1	1	13291	
0	5977	6	1	2	13282	1944	
0	5978	5	1	1	13283	
0	5979	6	1	2	13274	1945	
0	5980	5	1	1	13275	
0	5981	7	8	2	12824	13589	
0	5989	6	1	2	13186	1946	
0	5990	5	1	1	13187	
0	5991	6	4	2	5283	5284	
0	5996	6	3	2	5285	5286	
0	6000	6	2	2	5287	5288	
0	6003	6	5	2	5289	5290	
0	6009	6	4	2	5291	5292	
0	6014	6	3	2	5293	5294	
0	6018	6	2	2	5295	5296	
0	6021	6	1	2	5297	5298	
0	6022	6	1	2	5299	5300	
0	6023	5	1	1	13383	
0	6024	6	1	2	13384	4629	
0	6025	5	1	1	13378	
0	6026	6	1	2	13379	4631	
0	6027	5	1	1	13373	
0	6028	6	1	2	13374	4633	
0	6029	5	1	1	13363	
0	6030	6	1	2	13364	4636	
0	6031	5	1	1	13358	
0	6032	5	1	1	13230	
0	6033	5	1	1	13353	
0	6034	5	1	1	13225	
0	6035	5	1	1	13348	
0	6036	5	1	1	13220	
0	6037	5	1	1	13368	
0	6038	6	1	2	13369	4642	
0	6039	5	1	1	13343	
0	6040	5	1	1	13215	
0	6041	6	5	2	5314	5315	
0	6047	6	4	2	5316	5317	
0	6052	6	3	2	5318	5319	
0	6056	6	2	2	5320	5321	
0	6059	6	1	2	5322	5323	
0	6060	6	1	2	13336	1968	
0	6061	5	1	1	13337	
0	6062	6	1	2	13328	1969	
0	6063	5	1	1	13329	
0	6064	6	1	2	13320	1970	
0	6065	5	1	1	13321	
0	6066	6	1	2	13312	1971	
0	6067	5	1	1	13313	
0	6068	6	1	2	13302	1972	
0	6069	5	1	1	13303	
0	6070	6	1	2	13261	1973	
0	6071	5	1	1	13262	
0	6072	6	1	2	13253	1974	
0	6073	5	1	1	13254	
0	6074	6	1	2	13245	1975	
0	6075	5	1	1	13246	
0	6076	6	1	2	13237	1976	
0	6077	5	1	1	13238	
0	6078	5	1	1	13607	
0	6079	6	3	2	5363	4694	
0	6083	6	3	2	5364	5365	
0	6087	6	4	2	5366	5367	
0	6090	5	1	1	13239	
0	6091	6	1	2	13240	4699	
0	6092	5	1	1	13255	
0	6093	5	1	1	13247	
0	6094	5	1	1	13304	
0	6095	5	1	1	13263	
0	6096	5	1	1	13268	
0	6097	6	1	2	13269	4700	
0	6098	5	1	1	13284	
0	6099	5	1	1	13276	
0	6100	5	1	1	13178	
0	6101	5	1	1	13292	
0	6102	5	1	1	13609	
0	6103	6	1	2	13338	2015	
0	6104	5	1	1	13339	
0	6105	6	1	2	13330	2016	
0	6106	5	1	1	13331	
0	6107	6	1	2	13322	2017	
0	6108	5	1	1	13323	
0	6109	6	1	2	13305	2018	
0	6110	5	1	1	13306	
0	6111	6	1	2	13264	2019	
0	6112	5	1	1	13265	
0	6113	6	1	2	13256	2020	
0	6114	5	1	1	13257	
0	6115	6	1	2	13248	2021	
0	6116	5	1	1	13249	
0	6117	6	1	2	13314	2022	
0	6118	5	1	1	13315	
0	6119	6	1	2	13241	2023	
0	6120	5	1	1	13242	
0	6121	5	1	1	13216	
0	6122	6	1	2	13217	4743	
0	6123	5	1	1	13226	
0	6124	5	1	1	13221	
0	6125	6	1	2	13231	4744	
0	6126	5	1	1	13232	
0	6127	6	3	2	5425	4746	
0	6131	6	3	2	5426	5427	
0	6135	5	1	1	13148	
0	6136	6	1	2	13149	4749	
0	6137	6	3	2	5429	4751	
0	6141	6	3	2	5430	5431	
0	6145	6	4	2	5432	5433	
0	6148	5	1	1	13423	
0	6149	5	1	1	13168	
0	6150	5	1	1	13418	
0	6151	5	1	1	13163	
0	6152	5	1	1	13413	
0	6153	5	1	1	13158	
0	6154	5	1	1	13403	
0	6155	5	1	1	13150	
0	6156	5	1	1	13398	
0	6157	6	1	2	13399	4761	
0	6158	5	1	1	13393	
0	6159	6	1	2	13394	4763	
0	6160	5	1	1	13388	
0	6161	6	1	2	13389	4765	
0	6162	5	1	1	13408	
0	6163	5	1	1	13153	
0	6164	6	1	2	13298	4768	
0	6165	5	1	1	13299	
0	6166	6	3	2	5451	4776	
0	6170	6	3	2	5452	5453	
0	6174	6	4	2	5454	5455	
0	6177	6	3	2	5456	5457	
0	6181	5	1	1	13395	
0	6182	5	1	1	13390	
0	6183	5	1	1	13404	
0	6184	5	1	1	13400	
0	6185	5	1	1	13344	
0	6186	6	1	2	13345	4783	
0	6187	5	1	1	13354	
0	6188	5	1	1	13349	
0	6189	5	1	1	13365	
0	6190	5	1	1	13359	
0	6191	5	1	1	13595	
0	6192	6	1	2	13596	2230	
0	6193	5	1	1	13597	
0	6194	6	1	2	13598	2765	
0	6195	5	1	1	13043	
0	6196	6	2	2	5476	5477	
0	6199	6	2	2	5474	5475	
0	6202	5	1	1	13090	
0	6203	5	1	1	13110	
0	6213	5	1	1	13605	
0	6217	4	2	2	12825	13590	
0	6223	5	1	1	13324	
0	6224	5	1	1	13316	
0	6225	5	1	1	13340	
0	6226	5	1	1	13332	
0	6227	5	1	1	13196	
0	6228	5	1	1	13188	
0	6229	5	1	1	13212	
0	6230	5	1	1	13204	
0	6231	5	1	1	13611	
0	6235	5	1	1	13613	
0	6239	5	1	1	13159	
0	6240	5	1	1	13154	
0	6241	5	1	1	13169	
0	6242	5	1	1	13164	
0	6243	6	2	2	5573	5574	
0	6246	6	2	2	5571	5572	
0	6249	6	2	2	5586	5587	
0	6252	6	2	2	5584	5585	
0	6255	5	1	1	13414	
0	6256	5	1	1	13409	
0	6257	5	1	1	13424	
0	6258	5	1	1	13419	
0	6259	5	1	1	13375	
0	6260	5	1	1	13370	
0	6261	5	1	1	13385	
0	6262	5	1	1	13380	
0	6263	6	2	2	5604	5605	
0	6266	6	2	2	5602	5603	
0	6540	6	1	2	11863	5945	
0	6541	6	1	2	11854	5947	
0	6542	6	1	2	11847	5949	
0	6543	6	1	2	11834	5951	
0	6544	6	1	2	11825	5953	
0	6545	6	1	2	11816	5955	
0	6546	6	1	2	11809	5957	
0	6547	6	1	2	11800	5959	
0	6555	6	1	2	11864	5968	
0	6556	6	1	2	11855	5970	
0	6557	6	1	2	11848	5972	
0	6558	6	1	2	11826	5974	
0	6559	6	1	2	11817	5976	
0	6560	6	1	2	11810	5978	
0	6561	6	1	2	11801	5980	
0	6569	6	1	2	11835	5990	
0	6594	6	1	2	12861	6023	
0	6595	6	1	2	12854	6025	
0	6596	6	1	2	12849	6027	
0	6597	6	1	2	12836	6029	
0	6598	6	1	2	13233	6031	
0	6599	6	1	2	13360	6032	
0	6600	6	1	2	13227	6033	
0	6601	6	1	2	13355	6034	
0	6602	6	1	2	13222	6035	
0	6603	6	1	2	13350	6036	
0	6604	6	1	2	12844	6037	
0	6605	6	1	2	13218	6039	
0	6606	6	1	2	13346	6040	
0	6621	6	1	2	11939	6061	
0	6622	6	1	2	11932	6063	
0	6623	6	1	2	11925	6065	
0	6624	6	1	2	11918	6067	
0	6625	6	1	2	11907	6069	
0	6626	6	1	2	11897	6071	
0	6627	6	1	2	11890	6073	
0	6628	6	1	2	11883	6075	
0	6629	6	1	2	11876	6077	
0	6639	6	1	2	13438	6090	
0	6640	6	1	2	13250	6092	
0	6641	6	1	2	13258	6093	
0	6642	6	1	2	13266	6094	
0	6643	6	1	2	13307	6095	
0	6644	6	1	2	13440	6096	
0	6645	6	1	2	13277	6098	
0	6646	6	1	2	13285	6099	
0	6647	6	1	2	13293	6100	
0	6648	6	1	2	13179	6101	
0	6649	6	1	2	11940	6104	
0	6650	6	1	2	11933	6106	
0	6651	6	1	2	11926	6108	
0	6652	6	1	2	11908	6110	
0	6653	6	1	2	11898	6112	
0	6654	6	1	2	11891	6114	
0	6655	6	1	2	11884	6116	
0	6656	6	1	2	11919	6118	
0	6657	6	1	2	11877	6120	
0	6658	6	1	2	13444	6121	
0	6659	6	1	2	13223	6123	
0	6660	6	1	2	13228	6124	
0	6661	6	1	2	12837	6126	
0	6668	6	1	2	12743	6135	
0	6677	6	1	2	13170	6148	
0	6678	6	1	2	13425	6149	
0	6679	6	1	2	13165	6150	
0	6680	6	1	2	13420	6151	
0	6681	6	1	2	13160	6152	
0	6682	6	1	2	13415	6153	
0	6683	6	1	2	13151	6154	
0	6684	6	1	2	13405	6155	
0	6685	6	1	2	12744	6156	
0	6686	6	1	2	12735	6158	
0	6687	6	1	2	12728	6160	
0	6688	6	1	2	13155	6162	
0	6689	6	1	2	13410	6163	
0	6690	6	1	2	12830	6165	
0	6702	6	1	2	13391	6181	
0	6703	6	1	2	13396	6182	
0	6704	6	1	2	13401	6183	
0	6705	6	1	2	13406	6184	
0	6706	6	1	2	13460	6185	
0	6707	6	1	2	13351	6187	
0	6708	6	1	2	13356	6188	
0	6709	6	1	2	13361	6189	
0	6710	6	1	2	13366	6190	
0	6711	6	1	2	12250	6191	
0	6712	6	1	2	12217	6193	
0	6729	6	1	2	13317	6223	
0	6730	6	1	2	13325	6224	
0	6731	6	1	2	13333	6225	
0	6732	6	1	2	13341	6226	
0	6733	6	1	2	13189	6227	
0	6734	6	1	2	13197	6228	
0	6735	6	1	2	13205	6229	
0	6736	6	1	2	13213	6230	
0	6741	6	1	2	13156	6239	
0	6742	6	1	2	13161	6240	
0	6743	6	1	2	13166	6241	
0	6744	6	1	2	13171	6242	
0	6751	6	1	2	13411	6255	
0	6752	6	1	2	13416	6256	
0	6753	6	1	2	13421	6257	
0	6754	6	1	2	13426	6258	
0	6755	6	1	2	13371	6259	
0	6756	6	1	2	13376	6260	
0	6757	6	1	2	13381	6261	
0	6758	6	1	2	13386	6262	
0	6761	5	1	1	13895	
0	6762	7	3	5	13670	13656	13639	13624	13615	
0	6766	7	1	2	13616	13025	
0	6767	7	1	3	13625	13617	13028	
0	6768	7	1	4	13640	13618	13033	13626	
0	6769	7	1	5	13657	13641	13619	13044	13627	
0	6770	7	1	2	13628	13029	
0	6771	7	1	3	13642	13034	13629	
0	6772	7	1	4	13658	13643	13045	13630	
0	6773	7	1	4	13671	13644	13631	13659	
0	6774	7	1	2	13632	13030	
0	6775	7	1	3	13645	13035	13633	
0	6776	7	1	4	13660	13646	13046	13634	
0	6777	7	1	2	13647	13036	
0	6778	7	1	3	13661	13648	13047	
0	6779	7	1	3	13672	13649	13662	
0	6780	7	1	2	13650	13037	
0	6781	7	1	3	13663	13651	13048	
0	6782	7	1	2	13664	13049	
0	6783	7	1	2	13673	13665	
0	6784	7	2	5	13685	13716	13695	13678	13706	
0	6787	7	1	2	13679	13063	
0	6788	7	1	3	13686	13680	13065	
0	6789	7	1	4	13696	13681	13068	13687	
0	6790	7	1	5	13707	13697	13682	13072	13688	
0	6791	7	1	2	13689	13066	
0	6792	7	1	3	13698	13069	13690	
0	6793	7	1	4	13708	13699	13073	13691	
0	6794	7	1	2	13070	13700	
0	6795	7	1	3	13709	13701	13074	
0	6796	7	1	2	13710	13075	
0	6797	5	2	1	13723	
0	6800	5	2	1	13726	
0	6803	5	2	1	13733	
0	6806	5	2	1	13736	
0	6809	5	2	1	13743	
0	6812	5	2	1	13746	
0	6833	7	2	4	13846	13773	13761	13753	
0	6836	7	1	2	13754	13083	
0	6837	7	1	3	13762	13755	13086	
0	6838	7	1	4	13774	13756	13091	13763	
0	6839	7	1	2	13764	13087	
0	6840	7	1	3	13775	13092	13765	
0	6841	7	1	3	13847	13776	13766	
0	6842	7	1	2	13767	13088	
0	6843	7	1	3	13777	13093	13768	
0	6844	7	1	2	13778	13094	
0	6845	7	2	5	13853	13825	13808	13793	13784	
0	6848	7	1	2	13785	13096	
0	6849	7	1	3	13794	13786	13099	
0	6850	7	1	4	13809	13787	13104	13795	
0	6851	7	1	5	13826	13810	13788	13111	13796	
0	6852	7	1	2	13797	13100	
0	6853	7	1	3	13811	13105	13798	
0	6854	7	1	4	13827	13812	13112	13799	
0	6855	7	1	4	13854	13813	13800	13828	
0	6856	7	1	2	13801	13101	
0	6857	7	1	3	13814	13106	13802	
0	6858	7	1	4	13829	13815	13113	13803	
0	6859	7	1	2	13816	13107	
0	6860	7	1	3	13830	13817	13114	
0	6861	7	1	3	13855	13818	13831	
0	6862	7	1	2	13819	13108	
0	6863	7	1	3	13832	13820	13115	
0	6864	7	1	2	13833	13116	
0	6865	7	1	2	13848	13779	
0	6866	7	1	2	13856	13834	
0	6867	7	2	4	13869	13896	13881	13861	
0	6870	7	1	2	13862	13118	
0	6871	7	1	3	13870	13863	13121	
0	6872	7	1	4	13882	13864	13127	13871	
0	6873	7	1	2	13872	13122	
0	6874	7	1	3	13883	13128	13873	
0	6875	7	1	3	13897	13884	13874	
0	6876	7	1	2	13875	13123	
0	6877	7	1	3	13129	13885	13876	
0	6878	7	1	2	13886	13130	
0	6879	7	1	2	13898	13887	
0	6880	7	1	2	13888	13131	
0	6881	7	2	5	13907	13938	13917	13900	13928	
0	6884	7	1	2	13901	13133	
0	6885	7	1	3	13908	13902	13135	
0	6886	7	1	4	13918	13903	13138	13909	
0	6887	7	1	5	13929	13919	13904	13142	13910	
0	6888	7	1	2	13911	13136	
0	6889	7	1	3	13920	13139	13912	
0	6890	7	1	4	13930	13921	13143	13913	
0	6891	7	1	2	13140	13922	
0	6892	7	1	3	13931	13923	13144	
0	6893	7	1	2	13932	13145	
0	6894	6	8	2	5944	6540	
0	6901	6	12	2	5946	6541	
0	6912	6	12	2	5948	6542	
0	6923	6	5	2	5950	6543	
0	6929	6	7	2	5952	6544	
0	6936	6	10	2	5954	6545	
0	6946	6	11	2	5956	6546	
0	6957	6	10	2	5958	6547	
0	6967	6	1	2	13591	4575	
0	6968	5	1	1	13592	
0	6969	5	1	1	13481	
0	6970	6	8	2	5967	6555	
0	6977	6	12	2	5969	6556	
0	6988	6	11	2	5971	6557	
0	6998	6	9	2	5973	6558	
0	7006	6	15	2	5975	6559	
0	7020	6	17	2	5977	6560	
0	7036	6	14	2	5979	6561	
0	7049	6	7	2	5989	6569	
0	7055	6	1	2	13593	4610	
0	7056	5	1	1	13594	
0	7057	7	2	4	6021	13965	13962	13958	
0	7060	7	1	2	13959	3362	
0	7061	7	1	3	13963	13960	3363	
0	7062	7	1	4	13966	13961	3364	13964	
0	7063	7	1	5	6022	13979	13976	13972	13967	
0	7064	7	1	2	13968	3366	
0	7065	7	1	3	13973	13969	3367	
0	7066	7	1	4	13977	13970	3368	13974	
0	7067	7	1	5	13980	13978	13971	3369	13975	
0	7068	6	4	2	6594	6024	
0	7073	6	3	2	6595	6026	
0	7077	6	2	2	6596	6028	
0	7080	6	5	2	6597	6030	
0	7086	6	4	2	6598	6599	
0	7091	6	3	2	6600	6601	
0	7095	6	2	2	6602	6603	
0	7098	6	1	2	6604	6038	
0	7099	6	1	2	6605	6606	
0	7100	7	2	5	6059	13993	13990	13986	13981	
0	7103	7	1	2	13982	3371	
0	7104	7	1	3	13987	13983	3372	
0	7105	7	1	4	13991	13984	3373	13988	
0	7106	7	1	5	13994	13992	13985	3374	13989	
0	7107	6	8	2	6060	6621	
0	7114	6	12	2	6062	6622	
0	7125	6	12	2	6064	6623	
0	7136	6	5	2	6066	6624	
0	7142	6	7	2	6068	6625	
0	7149	6	10	2	6070	6626	
0	7159	6	11	2	6072	6627	
0	7170	6	10	2	6074	6628	
0	7180	6	7	2	6076	6629	
0	7187	5	1	1	13532	
0	7188	5	2	1	13995	
0	7191	5	2	1	13998	
0	7194	6	3	2	6639	6091	
0	7198	6	3	2	6640	6641	
0	7202	6	4	2	6642	6643	
0	7205	6	3	2	6644	6097	
0	7209	6	3	2	6645	6646	
0	7213	6	4	2	6647	6648	
0	7222	6	8	2	6103	6649	
0	7229	6	12	2	6105	6650	
0	7240	6	11	2	6107	6651	
0	7250	6	9	2	6109	6652	
0	7258	6	15	2	6111	6653	
0	7272	6	17	2	6113	6654	
0	7288	6	14	2	6115	6655	
0	7301	6	7	2	6117	6656	
0	7307	6	8	2	6119	6657	
0	7314	6	3	2	6658	6122	
0	7318	6	3	2	6659	6660	
0	7322	6	4	2	6125	6661	
0	7325	5	2	1	14005	
0	7328	5	2	1	14008	
0	7331	6	4	2	6668	6136	
0	7334	5	2	1	14011	
0	7337	5	2	1	14014	
0	7346	6	4	2	6677	6678	
0	7351	6	3	2	6679	6680	
0	7355	6	2	2	6681	6682	
0	7358	6	5	2	6683	6684	
0	7364	6	4	2	6685	6157	
0	7369	6	3	2	6686	6159	
0	7373	6	2	2	6687	6161	
0	7376	6	1	2	6688	6689	
0	7377	6	1	2	6164	6690	
0	7378	5	2	1	14021	
0	7381	5	2	1	14024	
0	7384	5	2	1	14031	
0	7387	6	3	2	6702	6703	
0	7391	6	4	2	6704	6705	
0	7394	6	3	2	6706	6186	
0	7398	6	3	2	6707	6708	
0	7402	6	4	2	6709	6710	
0	7441	6	2	2	6192	6711	
0	7444	6	2	2	6194	6712	
0	7477	5	1	1	14034	
0	7478	5	1	1	14036	
0	7551	5	1	1	13504	
0	7552	5	1	1	14038	
0	7556	5	1	1	14044	
0	7557	5	1	1	14046	
0	7558	5	1	1	14040	
0	7559	5	1	1	14042	
0	7560	6	2	2	6731	6732	
0	7563	6	2	2	6729	6730	
0	7566	6	2	2	6735	6736	
0	7569	6	2	2	6733	6734	
0	7572	5	1	1	13560	
0	7573	5	1	1	13580	
0	7574	6	2	2	6743	6744	
0	7577	6	2	2	6741	6742	
0	7580	5	1	1	14048	
0	7581	5	1	1	14050	
0	7582	6	2	2	6753	6754	
0	7585	6	2	2	6751	6752	
0	7588	6	2	2	6757	6758	
0	7591	6	2	2	6755	6756	
0	7609	3	3	5	3096	6766	6767	6768	6769	
0	7613	3	2	2	13038	6782	
0	7620	3	2	5	3136	6787	6788	6789	6790	
0	7649	3	1	4	3168	6836	6837	6838	
0	7650	3	2	2	13089	6844	
0	7655	3	3	5	3184	6848	6849	6850	6851	
0	7659	3	2	2	13109	6864	
0	7668	3	1	4	3210	6870	6871	6872	
0	7671	3	2	5	3228	6884	6885	6886	6887	
0	7744	6	1	2	12826	6968	
0	7822	6	1	2	12827	7056	
0	7825	3	1	4	3361	7060	7061	7062	
0	7826	3	1	5	3365	7064	7065	7066	7067	
0	7852	3	2	5	3370	7103	7104	7105	7106	
0	8114	3	2	4	13031	6777	6778	6779	
0	8117	3	2	5	13026	6770	6771	6772	6773	
0	8131	4	2	3	13032	6780	6781	
0	8134	4	2	4	13027	6774	6775	6776	
0	8144	6	1	2	14037	7477	
0	8145	6	1	2	14035	7478	
0	8146	3	2	4	13084	6839	6840	6841	
0	8156	4	2	3	13085	6842	6843	
0	8166	3	2	4	13102	6859	6860	6861	
0	8169	3	2	5	13097	6852	6853	6854	6855	
0	8183	4	2	3	13103	6862	6863	
0	8186	4	2	4	13098	6856	6857	6858	
0	8196	3	2	4	13119	6873	6874	6875	
0	8200	4	2	3	13120	6876	6877	
0	8204	3	2	3	13124	6878	6879	
0	8208	4	2	2	13125	6880	
0	8216	6	1	2	14047	7556	
0	8217	6	1	2	14045	7557	
0	8218	6	1	2	14043	7558	
0	8219	6	1	2	14041	7559	
0	8232	6	1	2	14051	7580	
0	8233	6	1	2	14049	7581	
0	8242	5	1	1	13939	
0	8243	5	1	1	13905	
0	8244	5	1	1	13914	
0	8245	5	1	1	13924	
0	8246	5	1	1	13933	
0	8247	5	1	1	13717	
0	8248	5	1	1	13683	
0	8249	5	1	1	13692	
0	8250	5	1	1	13702	
0	8251	5	1	1	13711	
0	8252	5	1	1	14304	
0	8253	5	1	1	14109	
0	8254	5	1	1	14052	
0	8260	5	1	1	13635	
0	8261	5	1	1	13636	
0	8262	7	4	2	13052	14053	
0	8269	7	4	2	13078	14055	
0	8274	5	1	1	13729	
0	8275	5	1	1	13730	
0	8276	5	1	1	13739	
0	8277	5	1	1	13740	
0	8278	5	1	1	13749	
0	8279	5	1	1	13750	
0	8280	7	1	3	13727	13724	13731	
0	8281	7	1	3	14059	14057	13732	
0	8282	7	1	3	13737	13734	13741	
0	8283	7	1	3	14063	14061	13742	
0	8284	7	1	3	13747	13744	13751	
0	8285	7	1	3	14067	14065	13752	
0	8288	5	1	1	14071	
0	8294	5	1	1	13769	
0	8295	5	1	1	13770	
0	8296	5	1	1	13804	
0	8297	5	1	1	13805	
0	8298	7	6	2	14069	14072	
0	8307	7	6	2	14073	14075	
0	8315	5	1	1	13865	
0	8317	5	1	1	13866	
0	8319	5	1	1	13877	
0	8321	5	1	1	13878	
0	8322	6	1	2	13889	4543	
0	8323	5	1	1	13890	
0	8324	6	1	2	13891	5943	
0	8325	5	1	1	13892	
0	8326	6	7	2	6967	7744	
0	8333	7	3	4	14085	14110	14097	14077	
0	8337	7	1	2	14078	13473	
0	8338	7	1	3	14086	14079	13476	
0	8339	7	1	4	14098	14080	13482	14087	
0	8340	7	1	2	14088	13477	
0	8341	7	1	3	14099	13483	14089	
0	8342	7	1	3	14111	14100	14090	
0	8343	7	1	2	14091	13478	
0	8344	7	1	3	13484	14101	14092	
0	8345	7	1	2	14102	13485	
0	8346	7	1	2	14112	14103	
0	8347	7	1	2	14104	13486	
0	8348	7	1	2	14114	13488	
0	8349	7	1	3	14121	14115	13490	
0	8350	7	1	4	14131	14116	13493	14122	
0	8351	7	1	5	14142	14132	14117	13945	14123	
0	8352	7	1	2	14124	13491	
0	8353	7	1	3	14133	13494	14125	
0	8354	7	1	4	14143	14134	13946	14126	
0	8355	7	1	2	13495	14135	
0	8356	7	1	3	14144	14136	13947	
0	8357	7	1	2	14145	13948	
0	8358	6	8	2	7055	7822	
0	8365	7	3	4	14238	14172	14160	14152	
0	8369	7	1	2	14153	13497	
0	8370	7	1	3	14161	14154	13500	
0	8371	7	1	4	14173	14155	13505	14162	
0	8372	7	1	2	14163	13501	
0	8373	7	1	3	14174	13506	14164	
0	8374	7	1	3	14239	14175	14165	
0	8375	7	1	2	14166	13502	
0	8376	7	1	3	14176	13507	14167	
0	8377	7	1	2	14177	13508	
0	8378	7	1	2	14183	13510	
0	8379	7	1	3	14192	14184	13513	
0	8380	7	1	4	14207	14185	13518	14193	
0	8381	7	1	5	14224	14208	14186	13950	14194	
0	8382	7	1	2	14195	13514	
0	8383	7	1	3	14209	13519	14196	
0	8384	7	1	4	14225	14210	13951	14197	
0	8385	7	1	2	14198	13515	
0	8386	7	1	3	14211	13520	14199	
0	8387	7	1	4	14226	14212	13952	14200	
0	8388	7	1	2	14213	13521	
0	8389	7	1	3	14227	14214	13953	
0	8390	7	1	2	14215	13522	
0	8391	7	1	3	14228	14216	13954	
0	8392	7	1	2	14229	13955	
0	8393	7	1	2	14240	14178	
0	8394	7	9	2	14245	7063	
0	8404	7	1	2	14246	7826	
0	8405	7	3	4	7098	14254	14251	14247	
0	8409	7	1	2	14248	4632	
0	8410	7	1	3	14252	14249	4634	
0	8411	7	1	4	14255	14250	4635	14253	
0	8412	7	2	5	7099	14268	14265	14261	14256	
0	8415	7	1	2	14257	4638	
0	8416	7	1	3	14262	14258	4639	
0	8417	7	1	4	14266	14259	4640	14263	
0	8418	7	1	5	14269	14267	14260	4641	14264	
0	8421	7	8	2	13295	14270	
0	8430	7	2	4	14280	14305	14292	14272	
0	8433	7	1	2	14273	13524	
0	8434	7	1	3	14281	14274	13527	
0	8435	7	1	4	14293	14275	13533	14282	
0	8436	7	1	2	14283	13528	
0	8437	7	1	3	14294	13534	14284	
0	8438	7	1	3	14306	14295	14285	
0	8439	7	1	2	14286	13529	
0	8440	7	1	3	13535	14296	14287	
0	8441	7	1	2	14297	13536	
0	8442	7	1	2	14307	14298	
0	8443	7	1	2	14299	13537	
0	8444	7	2	5	14316	14347	14326	14309	14337	
0	8447	7	1	2	14310	13539	
0	8448	7	1	3	14317	14311	13541	
0	8449	7	1	4	14327	14312	13544	14318	
0	8450	7	1	5	14338	14328	14313	13548	14319	
0	8451	7	1	2	14320	13542	
0	8452	7	1	3	14329	13545	14321	
0	8453	7	1	4	14339	14330	13549	14322	
0	8454	7	1	2	13546	14331	
0	8455	7	1	3	14340	14332	13550	
0	8456	7	1	2	14341	13551	
0	8457	5	2	1	14358	
0	8460	5	2	1	14361	
0	8463	5	2	1	14368	
0	8466	5	2	1	14371	
0	8469	5	1	1	14001	
0	8470	5	1	1	14002	
0	8483	7	1	3	13999	13996	14003	
0	8484	7	1	3	14356	14354	14004	
0	8485	7	2	4	14464	14398	14386	14378	
0	8488	7	1	2	14379	13553	
0	8489	7	1	3	14387	14380	13556	
0	8490	7	1	4	14399	14381	13561	14388	
0	8491	7	1	2	14389	13557	
0	8492	7	1	3	14400	13562	14390	
0	8493	7	1	3	14465	14401	14391	
0	8494	7	1	2	14392	13558	
0	8495	7	1	3	14402	13563	14393	
0	8496	7	1	2	14403	13564	
0	8497	7	2	5	14471	14450	14433	14418	14409	
0	8500	7	1	2	14410	13566	
0	8501	7	1	3	14419	14411	13569	
0	8502	7	1	4	14434	14412	13574	14420	
0	8503	7	1	5	14451	14435	14413	13581	14421	
0	8504	7	1	2	14422	13570	
0	8505	7	1	3	14436	13575	14423	
0	8506	7	1	4	14452	14437	13582	14424	
0	8507	7	1	4	14472	14438	14425	14453	
0	8508	7	1	2	14426	13571	
0	8509	7	1	3	14439	13576	14427	
0	8510	7	1	4	14454	14440	13583	14428	
0	8511	7	1	2	14441	13577	
0	8512	7	1	3	14455	14442	13584	
0	8513	7	1	3	14473	14443	14456	
0	8514	7	1	2	14444	13578	
0	8515	7	1	3	14457	14445	13585	
0	8516	7	1	2	14458	13586	
0	8517	7	1	2	14466	14404	
0	8518	7	1	2	14474	14459	
0	8519	5	2	1	14479	
0	8522	5	2	1	14482	
0	8537	5	1	1	14017	
0	8538	5	1	1	14018	
0	8539	7	1	3	14015	14012	14019	
0	8540	7	1	3	14499	14497	14020	
0	8541	7	3	4	7376	14508	14505	14501	
0	8545	7	1	2	14502	4757	
0	8546	7	1	3	14506	14503	4758	
0	8547	7	1	4	14509	14504	4759	14507	
0	8548	7	2	5	7377	14522	14519	14515	14510	
0	8551	7	1	2	14511	4762	
0	8552	7	1	3	14516	14512	4764	
0	8553	7	1	4	14520	14513	4766	14517	
0	8554	7	1	5	14523	14521	14514	4767	14518	
0	8555	5	2	1	14530	
0	8558	5	2	1	14537	
0	8561	5	2	1	14540	
0	8564	5	1	1	14027	
0	8565	5	1	1	14028	
0	8578	7	1	3	14025	14022	14029	
0	8579	7	1	3	14526	14524	14030	
0	8607	5	1	1	14547	
0	8608	6	1	2	14548	5469	
0	8609	5	1	1	14549	
0	8610	6	1	2	14550	4793	
0	8615	5	1	1	13674	
0	8616	5	1	1	13666	
0	8617	5	1	1	13620	
0	8618	5	1	1	13652	
0	8619	5	1	1	13653	
0	8624	5	1	1	13675	
0	8625	5	1	1	13667	
0	8626	5	1	1	13621	
0	8627	6	2	2	8144	8145	
0	8632	5	1	1	13849	
0	8633	5	1	1	13780	
0	8634	5	1	1	13757	
0	8637	5	1	1	13850	
0	8638	5	1	1	13781	
0	8639	5	1	1	13758	
0	8644	5	1	1	13857	
0	8645	5	1	1	13835	
0	8646	5	1	1	13789	
0	8647	5	1	1	13821	
0	8648	5	1	1	13822	
0	8653	5	1	1	13858	
0	8654	5	1	1	13836	
0	8655	5	1	1	13790	
0	8717	5	1	1	13956	
0	8727	6	2	2	8216	8217	
0	8730	6	2	2	8218	8219	
0	8733	5	1	1	14559	
0	8734	5	1	1	14561	
0	8753	5	1	1	14551	
0	8754	5	1	1	14553	
0	8755	5	1	1	14555	
0	8756	5	1	1	14557	
0	8811	6	2	2	8232	8233	
0	8814	5	1	1	14567	
0	8815	5	1	1	14569	
0	8816	5	1	1	14563	
0	8817	5	1	1	14565	
0	8818	7	1	2	14576	13079	
0	8840	7	1	2	13053	14571	
0	8857	5	3	1	14572	
0	8861	7	1	3	14058	13728	8274	
0	8862	7	1	3	13725	14060	8275	
0	8863	7	1	3	14062	13738	8276	
0	8864	7	1	3	13735	14064	8277	
0	8865	7	1	3	14066	13748	8278	
0	8866	7	1	3	13745	14068	8279	
0	8871	5	2	1	14580	
0	8874	7	1	2	14070	14581	
0	8878	7	1	2	14585	14074	
0	8879	5	1	1	11343	
0	8880	6	1	2	11344	8315	
0	8881	5	1	1	11348	
0	8882	6	1	2	11349	8317	
0	8883	5	1	1	11354	
0	8884	6	1	2	11355	8319	
0	8885	5	1	1	11359	
0	8886	6	1	2	11360	8321	
0	8887	6	1	2	13436	8323	
0	8888	6	1	2	13132	8325	
0	8898	3	3	4	4544	8337	8338	8339	
0	8902	3	2	5	4562	8348	8349	8350	8351	
0	8920	3	3	4	4576	8369	8370	8371	
0	8924	3	2	2	13503	8377	
0	8927	3	3	5	4592	8378	8379	8380	8381	
0	8931	3	2	2	13523	8392	
0	8943	3	3	2	7825	8404	
0	8950	3	3	4	4630	8409	8410	8411	
0	8956	3	2	5	4637	8415	8416	8417	8418	
0	8959	5	1	1	14587	
0	8960	7	1	2	13296	14588	
0	8963	3	1	4	4656	8433	8434	8435	
0	8966	3	2	5	4674	8447	8448	8449	8450	
0	8991	7	1	3	14355	14000	8469	
0	8992	7	1	3	13997	14357	8470	
0	8995	3	1	4	4701	8488	8489	8490	
0	8996	3	2	2	13559	8496	
0	9001	3	3	5	4717	8500	8501	8502	8503	
0	9005	3	2	2	13579	8516	
0	9024	7	1	3	14498	14016	8537	
0	9025	7	1	3	14013	14500	8538	
0	9029	3	3	4	4756	8545	8546	8547	
0	9035	3	2	5	4760	8551	8552	8553	8554	
0	9053	7	1	3	14525	14026	8564	
0	9054	7	1	3	14023	14527	8565	
0	9064	6	1	2	13472	8607	
0	9065	6	1	2	13428	8609	
0	9066	5	1	1	14589	
0	9067	6	1	2	14590	4795	
0	9068	3	2	2	14574	6783	
0	9071	5	1	1	14591	
0	9072	5	1	1	14593	
0	9073	6	1	2	14594	6195	
0	9074	5	2	1	14575	
0	9077	5	1	1	14595	
0	9079	3	2	2	14578	6865	
0	9082	5	1	1	14597	
0	9083	5	2	1	14579	
0	9086	5	1	1	14599	
0	9087	5	1	1	14601	
0	9088	6	1	2	14602	4813	
0	9089	3	2	2	14583	6866	
0	9092	5	1	1	14603	
0	9093	5	1	1	14605	
0	9094	6	1	2	14606	6203	
0	9095	5	2	1	14584	
0	9098	5	1	1	14607	
0	9099	3	2	4	13474	8340	8341	8342	
0	9103	4	2	3	13475	8343	8344	
0	9107	3	2	3	13479	8345	8346	
0	9111	4	2	2	13480	8347	
0	9117	3	2	4	13498	8372	8373	8374	
0	9127	4	2	3	13499	8375	8376	
0	9146	4	2	3	13516	8390	8391	
0	9149	4	2	4	13511	8385	8386	8387	
0	9159	6	1	2	14562	8733	
0	9160	6	1	2	14560	8734	
0	9161	3	2	4	13525	8436	8437	8438	
0	9165	4	2	3	13526	8439	8440	
0	9169	3	2	3	13530	8441	8442	
0	9173	4	2	2	13531	8443	
0	9179	6	1	2	14554	8753	
0	9180	6	1	2	14552	8754	
0	9181	6	1	2	14558	8755	
0	9182	6	1	2	14556	8756	
0	9183	3	2	4	13554	8491	8492	8493	
0	9193	4	2	3	13555	8494	8495	
0	9203	3	2	4	13572	8511	8512	8513	
0	9206	3	2	5	13567	8504	8505	8506	8507	
0	9220	4	2	3	13573	8514	8515	
0	9223	4	2	4	13568	8508	8509	8510	
0	9234	6	1	2	14570	8814	
0	9235	6	1	2	14568	8815	
0	9236	6	1	2	14566	8816	
0	9237	6	1	2	14564	8817	
0	9238	3	1	2	13081	8818	
0	9242	3	1	2	13055	8840	
0	9243	6	1	2	8324	8888	
0	9244	5	1	1	14348	
0	9245	5	1	1	14314	
0	9246	5	1	1	14323	
0	9247	5	1	1	14333	
0	9248	5	1	1	14342	
0	9249	5	1	1	14118	
0	9250	5	1	1	14127	
0	9251	5	1	1	14137	
0	9252	5	1	1	14146	
0	9256	4	1	2	8861	8280	
0	9257	4	1	2	8862	8281	
0	9258	4	1	2	8863	8282	
0	9259	4	1	2	8864	8283	
0	9260	4	1	2	8865	8284	
0	9261	4	1	2	8866	8285	
0	9262	5	1	1	11594	
0	9265	3	2	2	7649	8874	
0	9268	3	2	2	7668	8878	
0	9271	6	1	2	13867	8879	
0	9272	6	1	2	13868	8881	
0	9273	6	1	2	13879	8883	
0	9274	6	1	2	13880	8885	
0	9275	6	1	2	8322	8887	
0	9276	5	1	1	11520	
0	9280	7	2	5	14128	11511	14138	14119	14147	
0	9285	7	1	5	11572	11512	14139	14148	14129	
0	9286	7	1	4	11573	11513	14140	14149	
0	9287	7	1	3	11574	11514	14150	
0	9288	7	1	2	11575	11515	
0	9290	5	1	1	14081	
0	9292	5	1	1	14082	
0	9294	5	1	1	14093	
0	9296	5	1	1	14094	
0	9297	6	1	2	14105	5966	
0	9298	5	1	1	14106	
0	9299	6	1	2	14107	6969	
0	9300	5	1	1	14108	
0	9301	5	1	1	12017	
0	9307	7	3	5	12006	14230	14217	14201	14187	
0	9314	7	1	4	12007	14218	14202	14231	
0	9315	7	1	3	12008	14219	14232	
0	9318	7	1	2	12009	14233	
0	9319	5	1	1	14168	
0	9320	5	1	1	14169	
0	9321	5	1	1	14203	
0	9322	5	1	1	14204	
0	9323	5	1	1	11602	
0	9324	5	1	1	11604	
0	9326	5	1	1	12140	
0	9332	7	6	2	12141	12149	
0	9339	3	2	2	13469	8960	
0	9344	7	6	2	11527	11533	
0	9352	5	1	1	14276	
0	9354	5	1	1	14277	
0	9356	5	1	1	14288	
0	9358	5	1	1	14289	
0	9359	6	1	2	14300	6078	
0	9360	5	1	1	14301	
0	9361	6	1	2	14302	7187	
0	9362	5	1	1	14303	
0	9363	5	1	1	14364	
0	9364	5	1	1	14365	
0	9365	5	1	1	14374	
0	9366	5	1	1	14375	
0	9367	4	1	2	8991	8483	
0	9368	4	1	2	8992	8484	
0	9369	7	1	3	14362	14359	14366	
0	9370	7	1	3	11541	12233	14367	
0	9371	7	1	3	14372	14369	14376	
0	9372	7	1	3	11545	11543	14377	
0	9375	5	1	1	11555	
0	9381	5	1	1	14394	
0	9382	5	1	1	14395	
0	9383	5	1	1	14429	
0	9384	5	1	1	14430	
0	9385	7	6	2	11549	11556	
0	9392	5	1	1	14485	
0	9393	5	1	1	14486	
0	9394	5	1	1	14493	
0	9395	5	1	1	14494	
0	9396	7	1	3	14483	14480	14487	
0	9397	7	1	3	11559	11557	14488	
0	9398	7	1	3	14009	14006	14495	
0	9399	7	1	3	14491	14489	14496	
0	9400	4	1	2	9024	8539	
0	9401	4	1	2	9025	8540	
0	9402	5	1	1	11561	
0	9407	6	1	2	11564	11475	
0	9408	7	3	2	11562	11565	
0	9412	5	1	1	11636	
0	9413	5	1	1	14533	
0	9414	5	1	1	14534	
0	9415	5	1	1	14543	
0	9416	5	1	1	14544	
0	9417	4	1	2	9053	8578	
0	9418	4	1	2	9054	8579	
0	9419	7	1	3	14531	14032	14535	
0	9420	7	1	3	11566	14528	14536	
0	9421	7	1	3	14541	14538	14545	
0	9422	7	1	3	11588	11568	14546	
0	9426	6	2	2	9064	8608	
0	9429	6	2	2	9065	8610	
0	9432	6	1	2	13430	9066	
0	9435	6	1	2	13050	9072	
0	9442	6	1	2	13434	9087	
0	9445	6	1	2	13117	9093	
0	9454	5	1	1	14241	
0	9455	5	1	1	14179	
0	9456	5	1	1	14156	
0	9459	5	1	1	14242	
0	9460	5	1	1	14180	
0	9461	5	1	1	14157	
0	9465	5	1	1	14234	
0	9466	5	1	1	14188	
0	9467	5	1	1	14220	
0	9468	5	1	1	14221	
0	9476	5	1	1	14235	
0	9477	5	1	1	14189	
0	9478	6	2	2	9159	9160	
0	9485	6	2	2	9179	9180	
0	9488	6	2	2	9181	9182	
0	9493	5	1	1	14467	
0	9494	5	1	1	14405	
0	9495	5	1	1	14382	
0	9498	5	1	1	14468	
0	9499	5	1	1	14406	
0	9500	5	1	1	14383	
0	9505	5	1	1	14475	
0	9506	5	1	1	14460	
0	9507	5	1	1	14414	
0	9508	5	1	1	14446	
0	9509	5	1	1	14447	
0	9514	5	1	1	14476	
0	9515	5	1	1	14461	
0	9516	5	1	1	14415	
0	9517	6	2	2	9234	9235	
0	9520	6	2	2	9236	9237	
0	9526	7	1	2	11787	12154	
0	9531	7	1	2	11788	12155	
0	9539	6	1	2	9271	8880	
0	9540	6	1	2	9273	8884	
0	9541	5	1	1	9275	
0	9543	7	2	2	11690	8254	
0	9551	7	2	2	11700	8288	
0	9555	6	1	2	9272	8882	
0	9556	6	1	2	9274	8886	
0	9557	5	1	1	11722	
0	9560	7	1	2	11733	11521	
0	9561	5	1	1	11953	
0	9562	6	1	2	11954	9290	
0	9563	5	1	1	11955	
0	9564	6	1	2	11956	9292	
0	9565	5	1	1	11957	
0	9566	6	1	2	11958	9294	
0	9567	5	1	1	11959	
0	9568	6	1	2	11960	9296	
0	9569	6	1	2	13604	9298	
0	9570	6	1	2	13487	9300	
0	9571	5	1	1	11756	
0	9575	5	3	1	11770	
0	9579	7	1	2	12018	11771	
0	9581	5	1	1	11792	
0	9582	5	1	1	11802	
0	9585	7	1	2	12142	11803	
0	9591	7	1	2	11818	11528	
0	9592	5	1	1	11977	
0	9593	6	1	2	11978	9352	
0	9594	5	1	1	11979	
0	9595	6	1	2	11980	9354	
0	9596	5	1	1	11981	
0	9597	6	1	2	11982	9356	
0	9598	5	1	1	11983	
0	9599	6	1	2	11984	9358	
0	9600	6	1	2	13608	9360	
0	9601	6	1	2	13538	9362	
0	9602	7	1	3	12234	14363	9363	
0	9603	7	1	3	14360	11542	9364	
0	9604	7	1	3	11544	14373	9365	
0	9605	7	1	3	14370	11546	9366	
0	9608	5	2	1	11865	
0	9611	7	1	2	11550	11866	
0	9612	7	1	3	11558	14484	9392	
0	9613	7	1	3	14481	11560	9393	
0	9614	7	1	3	14490	14010	9394	
0	9615	7	1	3	14007	14492	9395	
0	9616	5	1	1	11899	
0	9617	5	1	1	11909	
0	9618	7	1	2	11563	11910	
0	9621	7	1	3	14529	14532	9413	
0	9622	7	1	3	14033	11567	9414	
0	9623	7	1	3	11569	14542	9415	
0	9624	7	1	3	14539	11589	9416	
0	9626	3	2	5	13489	8352	8353	8354	9285	
0	9629	3	2	4	13492	8355	8356	9286	
0	9632	3	2	3	13496	8357	9287	
0	9635	3	2	2	13949	9288	
0	9642	6	2	2	9067	9432	
0	9645	5	1	1	11941	
0	9646	6	2	2	9073	9435	
0	9649	5	1	1	11943	
0	9650	6	2	2	9257	9256	
0	9653	6	2	2	9259	9258	
0	9656	6	2	2	9261	9260	
0	9659	5	1	1	11945	
0	9660	6	1	2	11946	4809	
0	9661	5	1	1	11947	
0	9662	6	1	2	11948	6202	
0	9663	6	2	2	9088	9442	
0	9666	5	1	1	11949	
0	9667	6	2	2	9094	9445	
0	9670	5	1	1	11951	
0	9671	3	2	2	11759	8393	
0	9674	5	1	1	11961	
0	9675	5	2	1	11760	
0	9678	5	1	1	11963	
0	9679	3	2	4	13517	8388	8389	9315	
0	9682	3	2	2	11773	9318	
0	9685	3	2	5	13512	8382	8383	8384	9314	
0	9690	5	1	1	11965	
0	9691	6	1	2	11966	8717	
0	9692	5	2	1	11774	
0	9695	5	1	1	11975	
0	9698	6	2	2	9401	9400	
0	9702	6	2	2	9368	9367	
0	9707	3	2	2	11856	8517	
0	9710	5	1	1	11985	
0	9711	5	2	1	11857	
0	9714	5	1	1	11987	
0	9715	5	1	1	11989	
0	9716	6	1	2	11990	6235	
0	9717	3	2	2	11868	8518	
0	9720	5	1	1	11991	
0	9721	5	1	1	11996	
0	9722	6	1	2	11997	7573	
0	9723	5	2	1	11869	
0	9726	5	1	1	11998	
0	9727	6	2	2	9418	9417	
0	9732	7	1	2	12002	11672	
0	9733	6	1	2	9581	9326	
0	9734	7	1	5	11476	12110	12020	12123	12156	
0	9735	7	1	5	11477	12111	12021	12124	12157	
0	9736	7	1	2	12000	11632	
0	9737	5	1	1	9555	
0	9738	5	1	1	9556	
0	9739	6	1	2	9361	9601	
0	9740	6	1	2	11516	1115	
0	9741	5	1	1	11517	
0	9742	6	1	2	9299	9570	
0	9754	7	3	2	11522	12004	
0	9758	3	3	2	11723	9560	
0	9762	6	1	2	14083	9561	
0	9763	6	1	2	14084	9563	
0	9764	6	1	2	14095	9565	
0	9765	6	1	2	14096	9567	
0	9766	6	1	2	9297	9569	
0	9767	7	1	2	12005	11576	
0	9768	6	1	2	9557	9276	
0	9769	5	1	1	12014	
0	9773	6	1	2	12015	11577	
0	9774	6	1	2	9571	9301	
0	9775	7	3	2	12019	12016	
0	9779	3	3	2	11757	9579	
0	9784	5	1	1	12132	
0	9785	6	1	2	9616	9402	
0	9786	3	3	2	11793	9585	
0	9790	7	1	4	11478	12112	12022	12125	
0	9791	3	3	2	8963	9591	
0	9795	6	1	2	14278	9592	
0	9796	6	1	2	14279	9594	
0	9797	6	1	2	14290	9596	
0	9798	6	1	2	14291	9598	
0	9799	6	1	2	9359	9600	
0	9800	4	1	2	9602	9369	
0	9801	4	1	2	9603	9370	
0	9802	4	1	2	9604	9371	
0	9803	4	1	2	9605	9372	
0	9805	5	1	1	12134	
0	9806	5	1	1	12136	
0	9809	3	3	2	8995	9611	
0	9813	4	1	2	9612	9396	
0	9814	4	1	2	9613	9397	
0	9815	4	1	2	9614	9398	
0	9816	4	1	2	9615	9399	
0	9817	7	2	2	9617	9407	
0	9820	3	3	2	11900	9618	
0	9825	5	1	1	12138	
0	9826	5	1	1	12143	
0	9827	4	1	2	9621	9419	
0	9828	4	1	2	9622	9420	
0	9829	4	1	2	9623	9421	
0	9830	4	1	2	9624	9422	
0	9835	5	1	1	12119	
0	9836	6	1	2	12120	4789	
0	9837	5	1	1	12121	
0	9838	6	1	2	12122	4794	
0	9846	6	1	2	13432	9659	
0	9847	6	1	2	13095	9661	
0	9862	5	1	1	12010	
0	9863	6	1	2	13957	9690	
0	9866	5	1	1	12011	
0	9873	6	1	2	13614	9715	
0	9876	6	1	2	13587	9721	
0	9890	6	1	2	9795	9593	
0	9891	6	1	2	9797	9597	
0	9892	5	1	1	9799	
0	9893	6	1	2	11578	9741	
0	9894	6	1	2	9762	9562	
0	9895	6	1	2	9764	9566	
0	9896	5	1	1	9766	
0	9897	5	1	1	12164	
0	9898	6	1	2	12165	9249	
0	9899	5	1	1	12166	
0	9900	6	1	2	12167	9250	
0	9901	5	1	1	12168	
0	9902	6	1	2	12169	9251	
0	9903	5	1	1	12170	
0	9904	6	1	2	12171	9252	
0	9905	5	1	1	12145	
0	9906	5	1	1	12176	
0	9907	6	1	2	12177	5769	
0	9908	5	1	1	12178	
0	9909	6	1	2	12179	5770	
0	9910	5	1	1	12180	
0	9911	6	1	2	12181	9262	
0	9917	5	1	1	12147	
0	9923	6	1	2	9763	9564	
0	9924	6	1	2	9765	9568	
0	9925	3	6	2	11734	9767	
0	9932	7	2	2	12151	9773	
0	9935	7	2	2	12152	9769	
0	9938	5	1	1	12198	
0	9939	6	1	2	12199	9323	
0	9945	6	1	2	9796	9595	
0	9946	6	1	2	9798	9599	
0	9947	5	1	1	12200	
0	9948	6	1	2	12201	6102	
0	9949	7	2	2	12162	9375	
0	9953	5	1	1	12210	
0	9954	6	1	2	12211	9412	
0	9955	6	1	2	12653	9835	
0	9956	6	1	2	12654	9837	
0	9957	5	1	1	12172	
0	9958	6	1	2	12173	9645	
0	9959	5	1	1	12174	
0	9960	6	1	2	12175	9649	
0	9961	6	2	2	9660	9846	
0	9964	6	2	2	9662	9847	
0	9967	5	1	1	12182	
0	9968	6	1	2	12183	9666	
0	9969	5	1	1	12184	
0	9970	6	1	2	12185	9670	
0	9971	5	1	1	12186	
0	9972	6	1	2	12187	6213	
0	9973	5	1	1	12188	
0	9974	6	1	2	12189	7551	
0	9975	5	1	1	12190	
0	9976	6	1	2	12191	7552	
0	9977	5	1	1	12192	
0	9978	5	1	1	12194	
0	9979	6	2	2	9691	9863	
0	9982	5	1	1	12196	
0	9983	6	2	2	9814	9813	
0	9986	6	2	2	9816	9815	
0	9989	6	2	2	9801	9800	
0	9992	6	2	2	9803	9802	
0	9995	5	1	1	12202	
0	9996	6	1	2	12203	6231	
0	9997	5	1	1	12204	
0	9998	6	1	2	12205	7572	
0	9999	6	2	2	9716	9873	
0	10002	5	1	1	12206	
0	10003	6	2	2	9722	9876	
0	10006	5	1	1	12208	
0	10007	6	2	2	9830	9829	
0	10010	6	2	2	9828	9827	
0	10013	7	1	3	12238	11491	11673	
0	10014	7	1	4	12224	12028	11492	11674	
0	10015	7	1	5	11579	12221	12029	11493	11675	
0	10016	7	1	3	12235	12126	12158	
0	10017	7	1	4	12246	12023	12127	12159	
0	10018	7	1	3	12236	12128	12160	
0	10019	7	1	4	12247	12024	12129	12161	
0	10020	7	1	3	12241	11836	11633	
0	10021	7	1	4	12230	12068	11837	11634	
0	10022	7	1	5	11580	12227	12069	11838	11635	
0	10023	5	1	1	9945	
0	10024	5	1	1	9946	
3	10025	6	0	2	9740	9893	
0	10026	5	1	1	9923	
0	10028	5	1	1	9924	
0	10032	6	1	2	14120	9897	
0	10033	6	1	2	14130	9899	
0	10034	6	1	2	14141	9901	
0	10035	6	1	2	14151	9903	
0	10036	6	1	2	13600	9906	
0	10037	6	1	2	13602	9908	
0	10038	6	1	2	11595	9910	
0	10039	7	1	2	12242	11839	
0	10040	7	1	3	12231	12070	11840	
0	10041	7	1	4	11581	12228	12071	11841	
0	10042	7	1	2	12232	12072	
0	10043	7	1	3	11582	12229	12073	
0	10050	6	1	2	11603	9938	
0	10053	5	1	1	12244	
0	10054	7	1	2	12245	11901	
0	10055	7	1	2	12237	12130	
0	10056	7	1	3	12248	12025	12131	
0	10057	7	1	2	12239	11494	
0	10058	7	1	3	12225	12030	11495	
0	10059	7	1	4	11583	12222	12031	11496	
0	10060	7	1	2	12226	12032	
0	10061	7	1	3	11584	12223	12033	
0	10062	6	1	2	13610	9947	
0	10067	6	1	2	11637	9953	
0	10070	6	2	2	9955	9836	
0	10073	6	2	2	9956	9838	
0	10076	6	1	2	11942	9957	
0	10077	6	1	2	11944	9959	
0	10082	6	1	2	11950	9967	
0	10083	6	1	2	11952	9969	
0	10084	6	1	2	13606	9971	
0	10085	6	1	2	13509	9973	
0	10086	6	1	2	14039	9975	
0	10093	6	1	2	13612	9995	
0	10094	6	1	2	13565	9997	
3	10101	3	0	5	9238	9732	10013	10014	10015	
3	10102	3	0	5	12026	9526	10016	10017	9734	
3	10103	3	0	5	12027	9531	10018	10019	9735	
3	10104	3	0	5	9242	9736	10020	10021	10022	
0	10105	7	1	2	12253	9894	
0	10106	7	1	2	12254	9895	
0	10107	7	1	2	12255	9896	
0	10108	7	1	2	12256	8253	
3	10109	6	0	2	10032	9898	
3	10110	6	0	2	10033	9900	
3	10111	6	0	2	10034	9902	
3	10112	6	0	2	10035	9904	
0	10113	6	1	2	10036	9907	
0	10114	6	1	2	10037	9909	
0	10115	6	1	2	10038	9911	
0	10116	3	5	4	12001	10039	10040	10041	
0	10119	3	4	3	12243	10042	10043	
0	10124	5	5	1	12257	
0	10130	7	1	2	9768	12258	
0	10131	5	1	1	12259	
0	10132	5	1	1	12261	
0	10133	7	1	2	12260	11758	
0	10134	6	1	2	10050	9939	
0	10135	5	1	1	12288	
0	10136	6	1	2	12289	9324	
0	10137	5	1	1	12290	
0	10138	6	1	2	12291	9784	
0	10139	7	1	2	9785	10053	
0	10140	3	1	4	11789	10055	10056	9790	
0	10141	3	7	4	12003	10057	10058	10059	
0	10148	3	7	3	12240	10060	10061	
0	10155	6	1	2	10062	9948	
0	10156	5	1	1	12292	
0	10157	6	1	2	12293	9805	
0	10158	5	1	1	12294	
0	10159	6	1	2	12295	9806	
0	10160	5	1	1	12263	
0	10161	6	1	2	10067	9954	
0	10162	5	1	1	12303	
0	10163	6	1	2	12304	9825	
0	10164	5	1	1	12305	
0	10165	6	1	2	12306	9826	
0	10170	6	2	2	10076	9958	
0	10173	6	2	2	10077	9960	
0	10176	5	1	1	12269	
0	10177	6	1	2	12270	9082	
0	10178	5	1	1	12271	
0	10179	6	1	2	12272	9086	
0	10180	6	2	2	10082	9968	
0	10183	6	2	2	10083	9970	
0	10186	6	2	2	9972	10084	
0	10189	6	2	2	9974	10085	
0	10192	6	2	2	9976	10086	
0	10195	5	1	1	12281	
0	10196	6	1	2	12282	9982	
0	10197	6	2	2	9996	10093	
0	10200	6	2	2	9998	10094	
0	10203	5	1	1	12301	
0	10204	6	1	2	12302	10002	
0	10205	5	1	1	13893	
0	10206	6	1	2	13894	10006	
0	10212	6	1	2	12317	4308	
0	10213	6	1	2	12319	4313	
0	10230	7	1	2	9774	10131	
0	10231	6	1	2	11605	10135	
0	10232	6	1	2	12133	10137	
0	10233	3	1	2	10139	10054	
0	10234	6	1	2	14271	10140	
0	10237	6	1	2	12135	10156	
0	10238	6	1	2	12137	10158	
0	10239	6	1	2	12139	10162	
0	10240	6	1	2	12144	10164	
0	10241	5	1	1	12318	
0	10242	5	1	1	12320	
0	10247	6	1	2	14598	10176	
0	10248	6	1	2	14600	10178	
0	10259	6	1	2	12197	10195	
0	10264	6	1	2	12207	10203	
0	10265	6	1	2	12209	10205	
0	10266	7	1	2	10026	11782	
0	10267	7	1	2	10028	11783	
0	10268	7	1	2	9742	11784	
0	10269	7	1	2	14113	11785	
0	10270	6	1	2	14054	12326	
0	10271	6	1	2	12463	10241	
0	10272	6	1	2	12464	10242	
0	10278	7	1	5	13839	13718	13703	13712	13693	
0	10279	7	1	4	13840	13719	13704	13713	
0	10280	7	1	3	13841	13720	13714	
0	10281	7	1	2	13842	13721	
0	10282	7	1	2	14056	13843	
0	10283	5	3	1	12265	
0	10287	7	1	5	12339	13940	13925	13934	13915	
0	10288	7	1	4	12340	13941	13926	13935	
0	10289	7	1	3	12341	13942	13936	
0	10290	7	1	2	12342	13943	
0	10291	7	1	2	14076	12343	
0	10292	7	1	2	11724	11786	
0	10293	6	1	2	10231	10136	
0	10294	6	1	2	10232	10138	
0	10295	6	1	2	12150	10233	
0	10296	7	2	2	8959	10234	
0	10299	6	1	2	10237	10157	
0	10300	6	1	2	10238	10159	
0	10301	3	4	2	10230	10133	
0	10306	6	1	2	10239	10163	
0	10307	6	1	2	10240	10165	
0	10314	5	1	1	12356	
0	10315	6	1	2	12357	9071	
0	10316	5	1	1	12358	
0	10317	6	1	2	12359	9077	
0	10318	6	2	2	10247	10177	
0	10321	6	2	2	10248	10179	
0	10324	5	1	1	12387	
0	10325	6	1	2	12388	9092	
0	10326	5	1	1	12365	
0	10327	6	1	2	12366	9098	
0	10328	5	1	1	12367	
0	10329	6	1	2	12368	9674	
0	10330	5	1	1	12369	
0	10331	6	1	2	12370	9678	
0	10332	5	1	1	12371	
0	10333	6	1	2	12372	9977	
0	10334	6	2	2	10259	10196	
0	10337	5	1	1	12373	
0	10338	6	1	2	12374	9710	
0	10339	5	1	1	12375	
0	10340	6	1	2	12376	9714	
0	10341	6	2	2	10264	10204	
0	10344	6	2	2	10265	10206	
3	10350	3	0	2	10266	10105	
3	10351	3	0	2	10267	10106	
3	10352	3	0	2	10268	10107	
3	10353	3	0	2	10269	10108	
0	10354	7	2	2	11691	10270	
0	10357	6	2	2	10271	10212	
0	10360	6	2	2	10272	10213	
0	10367	3	4	2	14577	10282	
0	10375	3	5	2	14586	10291	
0	10381	3	7	2	10292	10130	
0	10388	7	2	4	10114	10134	10293	10294	
0	10391	7	2	2	9582	10295	
0	10399	7	2	4	10113	10115	10299	10300	
0	10402	7	2	4	10155	10161	10306	10307	
0	10406	3	2	5	13134	6888	6889	6890	10287	
0	10409	3	2	4	13137	6891	6892	10288	
0	10412	3	2	3	13141	6893	10289	
0	10415	3	2	2	13146	10290	
0	10419	3	2	5	13064	6791	6792	6793	10278	
0	10422	3	2	4	13067	6794	6795	10279	
0	10425	3	2	3	13071	6796	10280	
0	10428	3	2	2	13076	10281	
0	10431	6	1	2	14592	10314	
0	10432	6	1	2	14596	10316	
0	10437	6	1	2	14604	10324	
0	10438	6	1	2	14608	10326	
0	10439	6	1	2	11962	10328	
0	10440	6	1	2	11964	10330	
0	10441	6	1	2	12193	10332	
0	10444	6	1	2	11986	10337	
0	10445	6	1	2	11988	10339	
0	10450	5	1	1	12392	
0	10451	7	1	2	12393	13470	
0	10455	5	1	1	12344	
0	10456	6	1	2	12345	8242	
0	10465	5	1	1	13844	
0	10466	6	1	2	13845	8247	
0	10479	5	3	1	12327	
0	10497	5	3	1	12394	
0	10509	6	2	2	10431	10315	
0	10512	6	2	2	10432	10317	
0	10515	5	1	1	12398	
0	10516	6	1	2	12399	8632	
0	10517	5	1	1	12400	
0	10518	6	1	2	12401	8637	
0	10519	6	2	2	10437	10325	
0	10522	6	2	2	10438	10327	
0	10525	6	2	2	10439	10329	
0	10528	6	2	2	10440	10331	
0	10531	6	2	2	10441	10333	
0	10534	5	1	1	12402	
0	10535	6	1	2	12403	9695	
0	10536	6	2	2	10444	10338	
0	10539	6	2	2	10445	10340	
0	10542	5	1	1	12404	
0	10543	6	1	2	12405	9720	
0	10544	5	1	1	12406	
0	10545	6	1	2	12407	9726	
0	10546	7	1	2	5631	10450	
0	10547	5	1	1	12432	
0	10548	7	1	2	12433	11794	
0	10549	7	1	2	5165	12414	
0	10550	5	1	1	12408	
0	10551	7	1	2	12409	13056	
0	10552	6	1	2	13944	10455	
0	10553	7	1	2	12418	9539	
0	10554	7	1	2	12419	9540	
0	10555	7	1	2	12420	9541	
0	10556	7	1	2	12421	6761	
0	10557	5	1	1	12438	
0	10558	6	1	2	12439	8243	
0	10559	5	1	1	12440	
0	10560	6	1	2	12441	8244	
0	10561	5	1	1	12442	
0	10562	6	1	2	12443	8245	
0	10563	5	1	1	12444	
0	10564	6	1	2	12445	8246	
0	10565	6	1	2	13722	10465	
0	10566	5	1	1	12446	
0	10567	6	1	2	12447	8248	
0	10568	5	1	1	12448	
0	10569	6	1	2	12449	8249	
0	10570	5	1	1	12450	
0	10571	6	1	2	12451	8250	
0	10572	5	1	1	12452	
0	10573	6	1	2	12453	8251	
3	10574	5	0	1	12434	
3	10575	5	0	1	12436	
3	10576	5	0	1	12430	
0	10577	7	1	3	12435	12437	12431	
0	10581	7	1	3	12412	12146	12328	
0	10582	7	1	3	12410	9905	12329	
0	10583	5	3	1	12415	
0	10587	7	1	2	12416	5735	
0	10588	7	1	2	12417	3135	
0	10589	5	4	1	12422	
0	10594	7	1	5	12423	14349	14334	14343	14324	
0	10595	7	1	4	12424	14350	14335	14344	
0	10596	7	1	3	12425	14351	14345	
0	10597	7	1	2	12426	14352	
0	10598	7	1	2	11534	12427	
0	10609	6	1	2	13851	10515	
0	10610	6	1	2	13852	10517	
0	10621	6	1	2	11976	10534	
0	10626	6	1	2	11992	10542	
0	10627	6	1	2	11999	10544	
3	10628	3	0	2	10546	10451	
0	10629	7	1	2	9733	10547	
0	10631	7	1	2	5166	10550	
3	10632	6	0	2	10552	10456	
0	10637	6	1	2	13906	10557	
0	10638	6	1	2	13916	10559	
0	10639	6	1	2	13927	10561	
0	10640	6	1	2	13937	10563	
3	10641	6	0	2	10565	10466	
0	10642	6	1	2	13684	10566	
0	10643	6	1	2	13694	10568	
0	10644	6	1	2	13705	10570	
0	10645	6	1	2	13715	10572	
0	10647	7	1	3	886	887	10577	
0	10648	7	1	3	12413	11692	12476	
0	10649	7	1	3	12411	14573	12477	
0	10652	3	5	2	11819	10598	
0	10659	3	2	5	13540	8451	8452	8453	10594	
0	10662	3	2	4	13543	8454	8455	10595	
0	10665	3	2	3	13547	8456	10596	
0	10668	3	2	2	13552	10597	
0	10671	5	1	1	12497	
0	10672	6	1	2	12498	8615	
0	10673	5	1	1	12499	
0	10674	6	1	2	12500	8624	
0	10675	6	2	2	10609	10516	
0	10678	6	2	2	10610	10518	
0	10681	5	1	1	12506	
0	10682	6	1	2	12507	8644	
0	10683	5	1	1	13441	
0	10684	6	1	2	13442	8653	
0	10685	5	1	1	13445	
0	10686	6	1	2	13446	9454	
0	10687	5	1	1	13447	
0	10688	6	1	2	13448	9459	
0	10689	5	1	1	13449	
0	10690	6	1	2	13450	9978	
0	10691	6	2	2	10621	10535	
0	10694	5	1	1	13451	
0	10695	6	1	2	13452	9493	
0	10696	5	1	1	13453	
0	10697	6	1	2	13454	9498	
0	10698	6	2	2	10626	10543	
0	10701	6	2	2	10627	10545	
3	10704	3	0	2	10629	10548	
0	10705	7	1	2	13082	13461	
3	10706	3	0	2	10631	10551	
0	10707	7	1	2	9737	13464	
0	10708	7	1	2	9738	13465	
0	10709	7	1	2	9243	13466	
0	10710	7	1	2	13899	13467	
3	10711	6	0	2	10637	10558	
3	10712	6	0	2	10638	10560	
3	10713	6	0	2	10639	10562	
3	10714	6	0	2	10640	10564	
3	10715	6	0	2	10642	10567	
3	10716	6	0	2	10643	10569	
3	10717	6	0	2	10644	10571	
3	10718	6	0	2	10645	10573	
0	10719	5	1	1	12428	
0	10720	6	1	2	12429	9244	
3	10729	5	0	1	10647	
0	10730	7	1	2	5178	13462	
0	10731	7	1	2	12657	13463	
0	10737	6	1	2	13676	10671	
0	10738	6	1	2	13677	10673	
0	10739	3	2	4	10648	10649	10581	10582	
0	10746	6	1	2	13859	10681	
0	10747	6	1	2	13860	10683	
0	10748	6	1	2	14243	10685	
0	10749	6	1	2	14244	10687	
0	10750	6	1	2	12195	10689	
0	10753	6	1	2	14469	10694	
0	10754	6	1	2	14470	10696	
3	10759	3	0	2	10705	10549	
3	10760	3	0	2	10707	10553	
3	10761	3	0	2	10708	10554	
3	10762	3	0	2	10709	10555	
3	10763	3	0	2	10710	10556	
0	10764	6	1	2	14353	10719	
0	10765	7	1	2	12563	9890	
0	10766	7	1	2	12564	9891	
0	10767	7	1	2	12565	9892	
0	10768	7	1	2	12566	8252	
0	10769	5	1	1	12573	
0	10770	6	1	2	12574	9245	
0	10771	5	1	1	12580	
0	10772	6	1	2	12581	9246	
0	10773	5	1	1	12582	
0	10774	6	1	2	12583	9247	
0	10775	5	1	1	12589	
0	10776	6	1	2	12590	9248	
3	10778	3	0	2	10730	10587	
3	10781	3	0	2	10731	10588	
0	10784	5	4	1	12567	
0	10789	6	2	2	10737	10672	
0	10792	6	2	2	10738	10674	
0	10796	5	1	1	12604	
0	10797	6	1	2	12605	8633	
0	10798	5	1	1	12606	
0	10799	6	1	2	12607	8638	
0	10800	6	2	2	10746	10682	
0	10803	6	2	2	10747	10684	
0	10806	6	2	2	10748	10686	
0	10809	6	2	2	10749	10688	
0	10812	6	2	2	10750	10690	
0	10815	5	1	1	12626	
0	10816	6	1	2	12627	9866	
0	10817	6	2	2	10753	10695	
0	10820	6	2	2	10754	10697	
0	10823	5	1	1	12636	
0	10824	6	1	2	12637	9505	
0	10825	5	1	1	12646	
0	10826	6	1	2	12647	9514	
3	10827	6	0	2	10764	10720	
0	10832	6	1	2	14315	10769	
0	10833	6	1	2	14325	10771	
0	10834	6	1	2	14336	10773	
0	10835	6	1	2	14346	10775	
0	10836	5	1	1	12673	
0	10845	6	1	2	13782	10796	
0	10846	6	1	2	13783	10798	
0	10857	6	1	2	12012	10815	
0	10862	6	1	2	14477	10823	
0	10863	6	1	2	14478	10825	
0	10864	7	1	2	10023	12713	
0	10865	7	1	2	10024	12714	
0	10866	7	1	2	9739	12715	
0	10867	7	1	2	14308	12716	
3	10868	6	0	2	10832	10770	
3	10869	6	0	2	10833	10772	
3	10870	6	0	2	10834	10774	
3	10871	6	0	2	10835	10776	
0	10872	5	1	1	12717	
0	10873	6	1	2	12718	8616	
0	10874	5	1	1	12719	
0	10875	6	1	2	12720	8625	
0	10876	6	2	2	10845	10797	
0	10879	6	2	2	10846	10799	
0	10882	5	1	1	12729	
0	10883	6	1	2	12730	8645	
0	10884	5	1	1	12736	
0	10885	6	1	2	12737	8654	
0	10886	5	1	1	12738	
0	10887	6	1	2	12739	9455	
0	10888	5	1	1	12745	
0	10889	6	1	2	12746	9460	
0	10890	5	1	1	12756	
0	10891	6	1	2	12757	9862	
0	10892	6	2	2	10857	10816	
0	10895	5	1	1	12758	
0	10896	6	1	2	12759	9494	
0	10897	5	1	1	12768	
0	10898	6	1	2	12769	9499	
0	10899	6	2	2	10862	10824	
0	10902	6	2	2	10863	10826	
3	10905	3	0	2	10864	10765	
3	10906	3	0	2	10865	10766	
3	10907	3	0	2	10866	10767	
3	10908	3	0	2	10867	10768	
0	10909	6	1	2	13668	10872	
0	10910	6	1	2	13669	10874	
0	10915	6	1	2	13837	10882	
0	10916	6	1	2	13838	10884	
0	10917	6	1	2	14181	10886	
0	10918	6	1	2	14182	10888	
0	10919	6	1	2	12013	10890	
0	10922	6	1	2	14407	10895	
0	10923	6	1	2	14408	10897	
0	10928	6	2	2	10909	10873	
0	10931	6	2	2	10910	10875	
0	10934	5	1	1	12831	
0	10935	6	1	2	12832	8634	
0	10936	5	1	1	12838	
0	10937	6	1	2	12839	8639	
0	10938	6	2	2	10915	10883	
0	10941	6	2	2	10916	10885	
0	10944	6	2	2	10917	10887	
0	10947	6	2	2	10918	10889	
0	10950	6	2	2	10919	10891	
0	10953	5	1	1	12855	
0	10954	6	1	2	12856	9476	
0	10955	6	2	2	10922	10896	
0	10958	6	2	2	10923	10898	
0	10961	5	1	1	12862	
0	10962	6	1	2	12863	9506	
0	10963	5	1	1	12864	
0	10964	6	1	2	12865	9515	
0	10969	6	1	2	13759	10934	
0	10970	6	1	2	13760	10936	
0	10981	6	1	2	14236	10953	
0	10986	6	1	2	14462	10961	
0	10987	6	1	2	14463	10963	
0	10988	5	1	1	12876	
0	10989	6	1	2	12877	8617	
0	10990	5	1	1	12883	
0	10991	6	1	2	12884	8626	
0	10992	6	2	2	10969	10935	
0	10995	6	2	2	10970	10937	
0	10998	5	1	1	12895	
0	10999	6	1	2	12896	8646	
0	11000	5	1	1	12902	
0	11001	6	1	2	12903	8655	
0	11002	5	1	1	12904	
0	11003	6	1	2	12905	9456	
0	11004	5	1	1	12911	
0	11005	6	1	2	12912	9461	
0	11006	5	1	1	12918	
0	11007	6	1	2	12919	9465	
0	11008	6	2	2	10981	10954	
0	11011	5	1	1	12925	
0	11012	6	1	2	12926	9495	
0	11013	5	1	1	12929	
0	11014	6	1	2	12930	9500	
0	11015	6	2	2	10986	10962	
0	11018	6	2	2	10987	10964	
0	11023	6	1	2	13622	10988	
0	11024	6	1	2	13623	10990	
0	11027	6	1	2	13791	10998	
0	11028	6	1	2	13792	11000	
0	11029	6	1	2	14158	11002	
0	11030	6	1	2	14159	11004	
0	11031	6	1	2	14237	11006	
0	11034	6	1	2	14384	11011	
0	11035	6	1	2	14385	11013	
0	11040	5	1	1	12951	
0	11041	6	1	2	12952	8294	
0	11042	5	1	1	12953	
0	11043	6	1	2	12954	8295	
0	11044	6	2	2	11023	10989	
0	11047	6	2	2	11024	10991	
0	11050	6	2	2	11027	10999	
0	11053	6	2	2	11028	11001	
0	11056	6	2	2	11029	11003	
0	11059	6	2	2	11030	11005	
0	11062	6	2	2	11031	11007	
0	11065	5	1	1	12955	
0	11066	6	1	2	12956	9477	
0	11067	6	2	2	11034	11012	
0	11070	6	2	2	11035	11014	
0	11073	5	1	1	12957	
0	11074	6	1	2	12958	9507	
0	11075	5	1	1	12959	
0	11076	6	1	2	12960	9516	
0	11077	6	1	2	13771	11040	
0	11078	6	1	2	13772	11042	
0	11095	6	1	2	14190	11065	
0	11098	6	1	2	14416	11073	
0	11099	6	1	2	14417	11075	
0	11100	6	2	2	11077	11041	
0	11103	6	2	2	11078	11043	
0	11106	5	1	1	12969	
0	11107	6	1	2	12970	9319	
0	11108	5	1	1	12971	
0	11109	6	1	2	12972	9320	
0	11110	5	1	1	12975	
0	11111	6	1	2	12976	9381	
0	11112	5	1	1	12977	
0	11113	6	1	2	12978	9382	
0	11114	5	1	1	12961	
0	11115	6	1	2	12962	8618	
0	11116	5	1	1	12963	
0	11117	6	1	2	12964	8619	
0	11118	5	1	1	12965	
0	11119	6	1	2	12966	8647	
0	11120	5	1	1	12967	
0	11121	6	1	2	12968	8648	
0	11122	5	1	1	12973	
0	11123	6	1	2	12974	9466	
0	11124	6	2	2	11095	11066	
0	11127	6	2	2	11098	11074	
0	11130	6	2	2	11099	11076	
0	11137	6	1	2	14170	11106	
0	11138	6	1	2	14171	11108	
0	11139	6	1	2	14396	11110	
0	11140	6	1	2	14397	11112	
0	11141	6	1	2	13654	11114	
0	11142	6	1	2	13655	11116	
0	11143	6	1	2	13823	11118	
0	11144	6	1	2	13824	11120	
0	11145	6	1	2	14191	11122	
0	11152	7	1	3	12981	11701	12389	
0	11153	7	1	3	12979	14582	12390	
0	11154	7	1	3	12982	12148	12266	
0	11155	7	1	3	12980	9917	12267	
0	11156	6	2	2	11137	11107	
0	11159	6	2	2	11138	11109	
0	11162	6	2	2	11139	11111	
0	11165	6	2	2	11140	11113	
0	11168	6	2	2	11141	11115	
0	11171	6	2	2	11142	11117	
0	11174	6	2	2	11143	11119	
0	11177	6	2	2	11144	11121	
0	11180	6	2	2	11145	11123	
0	11183	5	1	1	12983	
0	11184	6	1	2	12984	9468	
0	11185	5	1	1	12985	
0	11186	6	1	2	12986	9508	
0	11187	5	1	1	12987	
0	11188	6	1	2	12988	9509	
0	11205	3	2	4	11152	11153	11154	11155	
0	11210	6	1	2	14222	11183	
0	11211	6	1	2	14448	11185	
0	11212	6	1	2	14449	11187	
0	11213	5	1	1	12997	
0	11214	6	1	2	12998	8260	
0	11215	5	1	1	12999	
0	11216	6	1	2	13000	8261	
0	11217	5	1	1	13001	
0	11218	6	1	2	13002	8296	
0	11219	5	1	1	13003	
0	11220	6	1	2	13004	8297	
0	11222	7	1	3	12991	12153	12113	
0	11223	7	1	3	12989	11772	12114	
0	11224	7	1	3	12992	12262	11585	
0	11225	7	1	3	12990	10132	11586	
0	11226	7	1	3	12995	12163	12489	
0	11227	7	1	3	12993	11867	12490	
0	11228	7	1	3	12996	12264	12395	
0	11229	7	1	3	12994	10160	12396	
0	11231	5	1	1	13005	
0	11232	6	1	2	13006	9467	
0	11233	6	2	2	11210	11184	
0	11236	6	2	2	11211	11186	
0	11239	6	2	2	11212	11188	
0	11242	6	1	2	13637	11213	
0	11243	6	1	2	13638	11215	
0	11244	6	1	2	13806	11217	
0	11245	6	1	2	13807	11219	
0	11246	5	1	1	13007	
0	11250	6	1	2	14223	11231	
0	11252	3	2	4	11222	11223	11224	11225	
0	11257	3	2	4	11226	11227	11228	11229	
0	11260	6	1	2	11242	11214	
0	11261	6	1	2	11243	11216	
0	11262	6	1	2	11244	11218	
0	11263	6	1	2	11245	11220	
0	11264	5	1	1	13009	
0	11265	6	1	2	13010	9322	
0	11267	5	1	1	13011	
0	11268	6	1	2	13012	9383	
0	11269	5	1	1	13013	
0	11270	6	1	2	13014	9384	
0	11272	6	2	2	11250	11232	
0	11277	5	1	1	11261	
0	11278	7	1	2	12330	11260	
0	11279	5	1	1	11263	
0	11280	7	1	2	12268	11262	
0	11282	6	1	2	14205	11264	
0	11283	5	1	1	13015	
0	11284	6	1	2	14431	11267	
0	11285	6	1	2	14432	11269	
0	11286	5	1	1	13017	
0	11288	7	1	2	11277	12478	
0	11289	7	1	2	11279	12391	
0	11290	5	1	1	13023	
0	11291	6	1	2	13024	9321	
0	11292	6	1	2	11282	11265	
0	11293	6	1	2	11284	11268	
0	11294	6	1	2	11285	11270	
0	11295	6	1	2	14206	11290	
0	11296	5	1	1	11292	
0	11297	5	1	1	11294	
0	11298	7	1	2	12397	11293	
0	11299	3	2	2	11288	11278	
0	11302	3	2	2	11289	11280	
0	11307	6	1	2	11295	11291	
0	11308	7	1	2	11296	12115	
0	11309	7	1	2	11297	12491	
0	11312	6	1	2	13041	11246	
0	11313	6	1	2	13039	10836	
0	11314	5	1	1	13040	
0	11315	5	1	1	13042	
0	11316	7	1	2	11587	11307	
0	11317	3	2	2	11309	11298	
0	11320	6	1	2	13008	11315	
0	11321	6	1	2	12674	11314	
0	11323	3	2	2	11308	11316	
0	11327	6	1	2	11312	11320	
0	11328	6	1	2	11313	11321	
0	11329	6	1	2	13057	11286	
0	11331	5	1	1	13058	
3	11333	5	0	1	11327	
3	11334	5	0	1	11328	
0	11335	6	1	2	13018	11331	
0	11336	6	1	2	13061	11283	
0	11337	5	1	1	13062	
0	11338	6	1	2	11329	11335	
0	11339	6	1	2	13016	11337	
3	11340	5	0	1	11338	
0	11341	6	1	2	11336	11339	
3	11342	5	0	1	11341	
2	11343	1	8196			
2	11344	1	8196			
2	11345	1	5			
2	11346	1	5			
2	11347	1	5			
2	11348	1	8200			
2	11349	1	8200			
2	11350	1	9			
2	11351	1	9			
2	11352	1	12			
2	11353	1	12			
2	11354	1	8204			
2	11355	1	8204			
2	11356	1	15			
2	11357	1	15			
2	11358	1	15			
2	11359	1	8208			
2	11360	1	8208			
2	11361	1	18			
2	11362	1	18			
2	11363	1	18			
2	11364	1	18			
2	11365	1	18			
2	11366	1	18			
2	11367	1	18			
2	11368	1	18			
2	11369	1	18			
2	11370	1	18			
2	11371	1	18			
2	11372	1	18			
2	11373	1	18			
2	11374	1	18			
2	11375	1	18			
2	11376	1	18			
2	11377	1	18			
2	11378	1	18			
2	11379	1	18			
2	11380	1	18			
2	11381	1	18			
2	11382	1	18			
2	11383	1	18			
2	11384	1	18			
2	11385	1	18			
2	11386	1	18			
2	11387	1	18			
2	11388	1	18			
2	11389	1	18			
2	11390	1	18			
2	11391	1	18			
2	11392	1	18			
2	11393	1	18			
2	11394	1	18			
2	11395	1	18			
2	11396	1	18			
2	11397	1	18			
2	11398	1	18			
2	11399	1	18			
2	11400	1	18			
2	11401	1	18			
2	11402	1	18			
2	11403	1	18			
2	11404	1	18			
2	11405	1	18			
2	11406	1	18			
2	11407	1	18			
2	11408	1	18			
2	11409	1	18			
2	11410	1	18			
2	11411	1	18			
2	11412	1	18			
2	11413	1	18			
2	11414	1	18			
2	11415	1	18			
2	11416	1	18			
2	11417	1	18			
2	11418	1	18			
2	11419	1	18			
2	11420	1	18			
2	11421	1	18			
2	11422	1	18			
2	11423	1	18			
2	11424	1	18			
2	11425	1	18			
2	11426	1	18			
2	11427	1	18			
2	11428	1	18			
2	11429	1	18			
2	11430	1	18			
2	11431	1	18			
2	11432	1	18			
2	11433	1	23			
2	11434	1	23			
2	11435	1	26			
2	11436	1	26			
2	11437	1	29			
2	11438	1	29			
2	11439	1	32			
2	11440	1	32			
2	11441	1	35			
2	11442	1	35			
2	11443	1	38			
2	11444	1	38			
2	11445	1	38			
2	11446	1	38			
2	11447	1	38			
2	11448	1	38			
2	11449	1	38			
2	11450	1	38			
2	11451	1	38			
2	11452	1	38			
2	11453	1	38			
2	11454	1	38			
2	11455	1	38			
2	11456	1	38			
2	11457	1	38			
2	11458	1	38			
2	11459	1	38			
2	11460	1	38			
2	11461	1	38			
2	11462	1	38			
2	11463	1	41			
2	11464	1	41			
2	11465	1	44			
2	11466	1	44			
2	11467	1	47			
2	11468	1	47			
2	11469	1	50			
2	11470	1	50			
2	11471	1	66			
2	11472	1	66			
2	11473	1	70			
2	11474	1	70			
2	11475	1	89			
2	11476	1	89			
2	11477	1	89			
2	11478	1	89			
2	11479	1	94			
2	11480	1	94			
2	11481	1	97			
2	11482	1	97			
2	11483	1	100			
2	11484	1	100			
2	11485	1	103			
2	11486	1	103			
2	11487	1	106			
2	11488	1	106			
2	11489	1	115			
2	11490	1	115			
2	11491	1	8307			
2	11492	1	8307			
2	11493	1	8307			
2	11494	1	8307			
2	11495	1	8307			
2	11496	1	8307			
2	11497	1	118			
2	11498	1	118			
2	11499	1	121			
2	11500	1	121			
2	11501	1	124			
2	11502	1	124			
2	11503	1	127			
2	11504	1	127			
2	11505	1	130			
2	11506	1	130			
2	11507	1	135			
2	11508	1	135			
2	11509	1	138			
2	11510	1	138			
2	11511	1	8326			
2	11512	1	8326			
2	11513	1	8326			
2	11514	1	8326			
2	11515	1	8326			
2	11516	1	8326			
2	11517	1	8326			
2	11518	1	141			
2	11519	1	141			
2	11520	1	8333			
2	11521	1	8333			
2	11522	1	8333			
2	11523	1	144			
2	11524	1	144			
2	11525	1	147			
2	11526	1	147			
2	11527	1	8430			
2	11528	1	8430			
2	11529	1	242			
2	11530	1	242			
2	11531	1	245			
2	11532	1	245			
2	11533	1	8444			
2	11534	1	8444			
2	11535	1	263			
2	11536	1	263			
2	11537	1	267			
2	11538	1	267			
2	11539	1	271			
2	11540	1	271			
2	11541	1	8460			
2	11542	1	8460			
2	11543	1	8463			
2	11544	1	8463			
2	11545	1	8466			
2	11546	1	8466			
2	11547	1	289			
2	11548	1	289			
2	11549	1	8485			
2	11550	1	8485			
2	11551	1	299			
2	11552	1	299			
2	11553	1	303			
2	11554	1	303			
2	11555	1	8497			
2	11556	1	8497			
2	11557	1	8519			
2	11558	1	8519			
2	11559	1	8522			
2	11560	1	8522			
2	11561	1	8541			
2	11562	1	8541			
2	11563	1	8541			
2	11564	1	8548			
2	11565	1	8548			
2	11566	1	8555			
2	11567	1	8555			
2	11568	1	8558			
2	11569	1	8558			
2	11570	1	367			
2	11571	1	367			
2	11572	1	367			
2	11573	1	367			
2	11574	1	367			
2	11575	1	367			
2	11576	1	367			
2	11577	1	367			
2	11578	1	367			
2	11579	1	367			
2	11580	1	367			
2	11581	1	367			
2	11582	1	367			
2	11583	1	367			
2	11584	1	367			
2	11585	1	367			
2	11586	1	367			
2	11587	1	367			
2	11588	1	8561			
2	11589	1	8561			
2	11590	1	382			
2	11591	1	382			
2	11592	1	382			
2	11593	1	382			
2	11594	1	8627			
2	11595	1	8627			
2	11596	1	469			
2	11597	1	469			
2	11598	1	494			
2	11599	1	494			
2	11600	1	528			
2	11601	1	528			
2	11602	1	8727			
2	11603	1	8727			
2	11604	1	8730			
2	11605	1	8730			
2	11606	1	575			
2	11607	1	575			
2	11608	1	578			
2	11609	1	578			
2	11610	1	593			
2	11611	1	593			
2	11612	1	596			
2	11613	1	596			
2	11614	1	599			
2	11615	1	599			
2	11616	1	599			
2	11617	1	599			
2	11618	1	599			
2	11619	1	599			
2	11620	1	604			
2	11621	1	604			
2	11622	1	604			
2	11623	1	604			
2	11624	1	604			
2	11625	1	604			
2	11626	1	609			
2	11627	1	609			
2	11628	1	609			
2	11629	1	609			
2	11630	1	609			
2	11631	1	609			
2	11632	1	8262			
2	11633	1	8262			
2	11634	1	8262			
2	11635	1	8262			
2	11636	1	8811			
2	11637	1	8811			
2	11638	1	628			
2	11639	1	628			
2	11640	1	628			
2	11641	1	628			
2	11642	1	628			
2	11643	1	628			
2	11644	1	628			
2	11645	1	628			
2	11646	1	628			
2	11647	1	628			
2	11648	1	628			
2	11649	1	628			
2	11650	1	628			
2	11651	1	632			
2	11652	1	632			
2	11653	1	632			
2	11654	1	632			
2	11655	1	632			
2	11656	1	632			
2	11657	1	632			
2	11658	1	632			
2	11659	1	632			
2	11660	1	632			
2	11661	1	632			
2	11662	1	632			
2	11663	1	632			
2	11664	1	644			
2	11665	1	644			
2	11666	1	644			
2	11667	1	644			
2	11668	1	644			
2	11669	1	644			
2	11670	1	644			
2	11671	1	644			
2	11672	1	8269			
2	11673	1	8269			
2	11674	1	8269			
2	11675	1	8269			
2	11676	1	651			
2	11677	1	651			
2	11678	1	651			
2	11679	1	651			
2	11680	1	651			
2	11681	1	651			
2	11682	1	651			
2	11683	1	660			
2	11684	1	660			
2	11685	1	660			
2	11686	1	660			
2	11687	1	660			
2	11688	1	660			
2	11689	1	660			
2	11690	1	8857			
2	11691	1	8857			
2	11692	1	8857			
2	11693	1	666			
2	11694	1	666			
2	11695	1	666			
2	11696	1	666			
2	11697	1	666			
2	11698	1	666			
2	11699	1	666			
2	11700	1	8871			
2	11701	1	8871			
2	11702	1	695			
2	11703	1	695			
2	11704	1	695			
2	11705	1	695			
2	11706	1	695			
2	11707	1	695			
2	11708	1	695			
2	11709	1	695			
2	11710	1	695			
2	11711	1	695			
2	11712	1	695			
2	11713	1	695			
2	11714	1	695			
2	11715	1	695			
2	11716	1	700			
2	11717	1	700			
2	11718	1	700			
2	11719	1	700			
2	11720	1	700			
2	11721	1	700			
2	11722	1	8898			
2	11723	1	8898			
2	11724	1	8898			
2	11725	1	708			
2	11726	1	708			
2	11727	1	708			
2	11728	1	708			
2	11729	1	708			
2	11730	1	708			
2	11731	1	708			
2	11732	1	708			
2	11733	1	8902			
2	11734	1	8902			
2	11735	1	715			
2	11736	1	715			
2	11737	1	715			
2	11738	1	715			
2	11739	1	715			
2	11740	1	715			
2	11741	1	715			
2	11742	1	721			
2	11743	1	721			
2	11744	1	721			
2	11745	1	721			
2	11746	1	721			
2	11747	1	721			
2	11748	1	721			
2	11749	1	727			
2	11750	1	727			
2	11751	1	727			
2	11752	1	727			
2	11753	1	727			
2	11754	1	727			
2	11755	1	727			
2	11756	1	8920			
2	11757	1	8920			
2	11758	1	8920			
2	11759	1	8924			
2	11760	1	8924			
2	11761	1	734			
2	11762	1	734			
2	11763	1	734			
2	11764	1	734			
2	11765	1	734			
2	11766	1	734			
2	11767	1	734			
2	11768	1	734			
2	11769	1	734			
2	11770	1	8927			
2	11771	1	8927			
2	11772	1	8927			
2	11773	1	8931			
2	11774	1	8931			
2	11775	1	742			
2	11776	1	742			
2	11777	1	742			
2	11778	1	742			
2	11779	1	742			
2	11780	1	742			
2	11781	1	742			
2	11782	1	10124			
2	11783	1	10124			
2	11784	1	10124			
2	11785	1	10124			
2	11786	1	10124			
2	11787	1	8943			
2	11788	1	8943			
2	11789	1	8943			
2	11790	1	759			
2	11791	1	759			
2	11792	1	8950			
2	11793	1	8950			
2	11794	1	8950			
2	11795	1	762			
2	11796	1	762			
2	11797	1	762			
2	11798	1	762			
2	11799	1	762			
2	11800	1	762			
2	11801	1	762			
2	11802	1	8956			
2	11803	1	8956			
2	11804	1	768			
2	11805	1	768			
2	11806	1	768			
2	11807	1	768			
2	11808	1	768			
2	11809	1	768			
2	11810	1	768			
2	11811	1	774			
2	11812	1	774			
2	11813	1	774			
2	11814	1	774			
2	11815	1	774			
2	11816	1	774			
2	11817	1	774			
2	11818	1	8966			
2	11819	1	8966			
2	11820	1	780			
2	11821	1	780			
2	11822	1	780			
2	11823	1	780			
2	11824	1	780			
2	11825	1	780			
2	11826	1	780			
2	11827	1	786			
2	11828	1	786			
2	11829	1	786			
2	11830	1	786			
2	11831	1	786			
2	11832	1	786			
2	11833	1	786			
2	11834	1	786			
2	11835	1	786			
2	11836	1	8298			
2	11837	1	8298			
2	11838	1	8298			
2	11839	1	8298			
2	11840	1	8298			
2	11841	1	8298			
2	11842	1	794			
2	11843	1	794			
2	11844	1	794			
2	11845	1	794			
2	11846	1	794			
2	11847	1	794			
2	11848	1	794			
2	11849	1	800			
2	11850	1	800			
2	11851	1	800			
2	11852	1	800			
2	11853	1	800			
2	11854	1	800			
2	11855	1	800			
2	11856	1	8996			
2	11857	1	8996			
2	11858	1	806			
2	11859	1	806			
2	11860	1	806			
2	11861	1	806			
2	11862	1	806			
2	11863	1	806			
2	11864	1	806			
2	11865	1	9001			
2	11866	1	9001			
2	11867	1	9001			
2	11868	1	9005			
2	11869	1	9005			
2	11870	1	814			
2	11871	1	814			
2	11872	1	814			
2	11873	1	814			
2	11874	1	814			
2	11875	1	814			
2	11876	1	814			
2	11877	1	814			
2	11878	1	821			
2	11879	1	821			
2	11880	1	821			
2	11881	1	821			
2	11882	1	821			
2	11883	1	821			
2	11884	1	821			
2	11885	1	827			
2	11886	1	827			
2	11887	1	827			
2	11888	1	827			
2	11889	1	827			
2	11890	1	827			
2	11891	1	827			
2	11892	1	833			
2	11893	1	833			
2	11894	1	833			
2	11895	1	833			
2	11896	1	833			
2	11897	1	833			
2	11898	1	833			
2	11899	1	9029			
2	11900	1	9029			
2	11901	1	9029			
2	11902	1	839			
2	11903	1	839			
2	11904	1	839			
2	11905	1	839			
2	11906	1	839			
2	11907	1	839			
2	11908	1	839			
2	11909	1	9035			
2	11910	1	9035			
2	11911	1	845			
2	11912	1	845			
2	11913	1	845			
2	11914	1	845			
2	11915	1	845			
2	11916	1	845			
2	11917	1	845			
2	11918	1	845			
2	11919	1	845			
2	11920	1	853			
2	11921	1	853			
2	11922	1	853			
2	11923	1	853			
2	11924	1	853			
2	11925	1	853			
2	11926	1	853			
2	11927	1	859			
2	11928	1	859			
2	11929	1	859			
2	11930	1	859			
2	11931	1	859			
2	11932	1	859			
2	11933	1	859			
2	11934	1	865			
2	11935	1	865			
2	11936	1	865			
2	11937	1	865			
2	11938	1	865			
2	11939	1	865			
2	11940	1	865			
2	11941	1	9068			
2	11942	1	9068			
2	11943	1	9074			
2	11944	1	9074			
2	11945	1	9079			
2	11946	1	9079			
2	11947	1	9083			
2	11948	1	9083			
2	11949	1	9089			
2	11950	1	9089			
2	11951	1	9095			
2	11952	1	9095			
2	11953	1	9099			
2	11954	1	9099			
2	11955	1	9103			
2	11956	1	9103			
2	11957	1	9107			
2	11958	1	9107			
2	11959	1	9111			
2	11960	1	9111			
2	11961	1	9117			
2	11962	1	9117			
2	11963	1	9127			
2	11964	1	9127			
2	11965	1	9146			
2	11966	1	9146			
2	11967	1	957			
2	11968	1	957			
2	11969	1	957			
2	11970	1	957			
2	11971	1	957			
2	11972	1	957			
2	11973	1	957			
2	11974	1	957			
2	11975	1	9149			
2	11976	1	9149			
2	11977	1	9161			
2	11978	1	9161			
2	11979	1	9165			
2	11980	1	9165			
2	11981	1	9169			
2	11982	1	9169			
2	11983	1	9173			
2	11984	1	9173			
2	11985	1	9183			
2	11986	1	9183			
2	11987	1	9193			
2	11988	1	9193			
2	11989	1	9203			
2	11990	1	9203			
2	11991	1	9206			
2	11992	1	9206			
2	11993	1	1029			
2	11994	1	1029			
2	11995	1	1029			
2	11996	1	9220			
2	11997	1	9220			
2	11998	1	9223			
2	11999	1	9223			
2	12000	1	9265			
2	12001	1	9265			
2	12002	1	9268			
2	12003	1	9268			
2	12004	1	9280			
2	12005	1	9280			
2	12006	1	8358			
2	12007	1	8358			
2	12008	1	8358			
2	12009	1	8358			
2	12010	1	8358			
2	12011	1	8358			
2	12012	1	8358			
2	12013	1	8358			
2	12014	1	9307			
2	12015	1	9307			
2	12016	1	9307			
2	12017	1	8365			
2	12018	1	8365			
2	12019	1	8365			
2	12020	1	9332			
2	12021	1	9332			
2	12022	1	9332			
2	12023	1	9332			
2	12024	1	9332			
2	12025	1	9332			
2	12026	1	9339			
2	12027	1	9339			
2	12028	1	9344			
2	12029	1	9344			
2	12030	1	9344			
2	12031	1	9344			
2	12032	1	9344			
2	12033	1	9344			
2	12034	1	1167			
2	12035	1	1167			
2	12036	1	1167			
2	12037	1	1167			
2	12038	1	1189			
2	12039	1	1189			
2	12040	1	1189			
2	12041	1	1189			
2	12042	1	1189			
2	12043	1	1189			
2	12044	1	1194			
2	12045	1	1194			
2	12046	1	1194			
2	12047	1	1194			
2	12048	1	1194			
2	12049	1	1194			
2	12050	1	1194			
2	12051	1	1194			
2	12052	1	1194			
2	12053	1	1194			
2	12054	1	1194			
2	12055	1	1194			
2	12056	1	1194			
2	12057	1	1194			
2	12058	1	1194			
2	12059	1	1194			
2	12060	1	1194			
2	12061	1	1194			
2	12062	1	1194			
2	12063	1	1194			
2	12064	1	1194			
2	12065	1	1194			
2	12066	1	1194			
2	12067	1	1194			
2	12068	1	9385			
2	12069	1	9385			
2	12070	1	9385			
2	12071	1	9385			
2	12072	1	9385			
2	12073	1	9385			
2	12074	1	1199			
2	12075	1	1199			
2	12076	1	1199			
2	12077	1	1199			
2	12078	1	1199			
2	12079	1	1199			
2	12080	1	1199			
2	12081	1	1199			
2	12082	1	1199			
2	12083	1	1199			
2	12084	1	1199			
2	12085	1	1199			
2	12086	1	1206			
2	12087	1	1206			
2	12088	1	1206			
2	12089	1	1206			
2	12090	1	1206			
2	12091	1	1206			
2	12092	1	1206			
2	12093	1	1206			
2	12094	1	1206			
2	12095	1	1206			
2	12096	1	1206			
2	12097	1	1206			
2	12098	1	1206			
2	12099	1	1206			
2	12100	1	1206			
2	12101	1	1206			
2	12102	1	1206			
2	12103	1	1206			
2	12104	1	1206			
2	12105	1	1206			
2	12106	1	1206			
2	12107	1	1206			
2	12108	1	1206			
2	12109	1	1206			
2	12110	1	9408			
2	12111	1	9408			
2	12112	1	9408			
2	12113	1	1218			
2	12114	1	1218			
2	12115	1	1218			
2	12116	1	1222			
2	12117	1	1222			
2	12118	1	1222			
2	12119	1	9426			
2	12120	1	9426			
2	12121	1	9429			
2	12122	1	9429			
2	12123	1	8394			
2	12124	1	8394			
2	12125	1	8394			
2	12126	1	8394			
2	12127	1	8394			
2	12128	1	8394			
2	12129	1	8394			
2	12130	1	8394			
2	12131	1	8394			
2	12132	1	9478			
2	12133	1	9478			
2	12134	1	9485			
2	12135	1	9485			
2	12136	1	9488			
2	12137	1	9488			
2	12138	1	9517			
2	12139	1	9517			
2	12140	1	8405			
2	12141	1	8405			
2	12142	1	8405			
2	12143	1	9520			
2	12144	1	9520			
2	12145	1	9543			
2	12146	1	9543			
2	12147	1	9551			
2	12148	1	9551			
2	12149	1	8412			
2	12150	1	8412			
2	12151	1	9575			
2	12152	1	9575			
2	12153	1	9575			
2	12154	1	8421			
2	12155	1	8421			
2	12156	1	8421			
2	12157	1	8421			
2	12158	1	8421			
2	12159	1	8421			
2	12160	1	8421			
2	12161	1	8421			
2	12162	1	9608			
2	12163	1	9608			
2	12164	1	9626			
2	12165	1	9626			
2	12166	1	9629			
2	12167	1	9629			
2	12168	1	9632			
2	12169	1	9632			
2	12170	1	9635			
2	12171	1	9635			
2	12172	1	9642			
2	12173	1	9642			
2	12174	1	9646			
2	12175	1	9646			
2	12176	1	9650			
2	12177	1	9650			
2	12178	1	9653			
2	12179	1	9653			
2	12180	1	9656			
2	12181	1	9656			
2	12182	1	9663			
2	12183	1	9663			
2	12184	1	9667			
2	12185	1	9667			
2	12186	1	9671			
2	12187	1	9671			
2	12188	1	9675			
2	12189	1	9675			
2	12190	1	9679			
2	12191	1	9679			
2	12192	1	9682			
2	12193	1	9682			
2	12194	1	9685			
2	12195	1	9685			
2	12196	1	9692			
2	12197	1	9692			
2	12198	1	9698			
2	12199	1	9698			
2	12200	1	9702			
2	12201	1	9702			
2	12202	1	9707			
2	12203	1	9707			
2	12204	1	9711			
2	12205	1	9711			
2	12206	1	9717			
2	12207	1	9717			
2	12208	1	9723			
2	12209	1	9723			
2	12210	1	9727			
2	12211	1	9727			
2	12212	1	1537			
2	12213	1	1537			
2	12214	1	1537			
2	12215	1	1537			
2	12216	1	1537			
2	12217	1	1537			
2	12218	1	1551			
2	12219	1	1551			
2	12220	1	1551			
2	12221	1	9754			
2	12222	1	9754			
2	12223	1	9754			
2	12224	1	9758			
2	12225	1	9758			
2	12226	1	9758			
2	12227	1	9775			
2	12228	1	9775			
2	12229	1	9775			
2	12230	1	9779			
2	12231	1	9779			
2	12232	1	9779			
2	12233	1	8457			
2	12234	1	8457			
2	12235	1	9786			
2	12236	1	9786			
2	12237	1	9786			
2	12238	1	9791			
2	12239	1	9791			
2	12240	1	9791			
2	12241	1	9809			
2	12242	1	9809			
2	12243	1	9809			
2	12244	1	9817			
2	12245	1	9817			
2	12246	1	9820			
2	12247	1	9820			
2	12248	1	9820			
2	12249	1	1708			
2	12250	1	1708			
2	12251	1	1721			
2	12252	1	1721			
2	12253	1	9925			
2	12254	1	9925			
2	12255	1	9925			
2	12256	1	9925			
2	12257	1	9925			
2	12258	1	9925			
2	12259	1	9932			
2	12260	1	9932			
2	12261	1	9935			
2	12262	1	9935			
2	12263	1	9949			
2	12264	1	9949			
2	12265	1	10119			
2	12266	1	10119			
2	12267	1	10119			
2	12268	1	10119			
2	12269	1	9961			
2	12270	1	9961			
2	12271	1	9964			
2	12272	1	9964			
2	12273	1	1783			
2	12274	1	1783			
2	12275	1	1783			
2	12276	1	1783			
2	12277	1	1783			
2	12278	1	1789			
2	12279	1	1789			
2	12280	1	1789			
2	12281	1	9979			
2	12282	1	9979			
2	12283	1	1799			
2	12284	1	1799			
2	12285	1	1799			
2	12286	1	1799			
2	12287	1	1799			
2	12288	1	9983			
2	12289	1	9983			
2	12290	1	9986			
2	12291	1	9986			
2	12292	1	9989			
2	12293	1	9989			
2	12294	1	9992			
2	12295	1	9992			
2	12296	1	1805			
2	12297	1	1805			
2	12298	1	1805			
2	12299	1	1805			
2	12300	1	1805			
2	12301	1	9999			
2	12302	1	9999			
2	12303	1	10007			
2	12304	1	10007			
2	12305	1	10010			
2	12306	1	10010			
2	12307	1	1845			
2	12308	1	1845			
2	12309	1	1845			
2	12310	1	1845			
2	12311	1	1845			
2	12312	1	1851			
2	12313	1	1851			
2	12314	1	1851			
2	12315	1	1851			
2	12316	1	1851			
2	12317	1	10070			
2	12318	1	10070			
2	12319	1	10073			
2	12320	1	10073			
2	12321	1	1913			
2	12322	1	1913			
2	12323	1	1913			
2	12324	1	1913			
2	12325	1	1913			
2	12326	1	10116			
2	12327	1	10116			
2	12328	1	10116			
2	12329	1	10116			
2	12330	1	10116			
2	12331	1	1947			
2	12332	1	1947			
2	12333	1	1947			
2	12334	1	1947			
2	12335	1	1947			
2	12336	1	1953			
2	12337	1	1953			
2	12338	1	1953			
2	12339	1	10148			
2	12340	1	10148			
2	12341	1	10148			
2	12342	1	10148			
2	12343	1	10148			
2	12344	1	10148			
2	12345	1	10148			
2	12346	1	1977			
2	12347	1	1977			
2	12348	1	1977			
2	12349	1	1977			
2	12350	1	1977			
2	12351	1	1983			
2	12352	1	1983			
2	12353	1	1983			
2	12354	1	1983			
2	12355	1	1983			
2	12356	1	10170			
2	12357	1	10170			
2	12358	1	10173			
2	12359	1	10173			
2	12360	1	1997			
2	12361	1	1997			
2	12362	1	1997			
2	12363	1	1997			
2	12364	1	1997			
2	12365	1	10183			
2	12366	1	10183			
2	12367	1	10186			
2	12368	1	10186			
2	12369	1	10189			
2	12370	1	10189			
2	12371	1	10192			
2	12372	1	10192			
2	12373	1	10197			
2	12374	1	10197			
2	12375	1	10200			
2	12376	1	10200			
2	12377	1	2052			
2	12378	1	2052			
2	12379	1	2052			
2	12380	1	2052			
2	12381	1	2052			
2	12382	1	2058			
2	12383	1	2058			
2	12384	1	2058			
2	12385	1	2058			
2	12386	1	2058			
2	12387	1	10180			
2	12388	1	10180			
2	12389	1	10283			
2	12390	1	10283			
2	12391	1	10283			
2	12392	1	10296			
2	12393	1	10296			
2	12394	1	10301			
2	12395	1	10301			
2	12396	1	10301			
2	12397	1	10301			
2	12398	1	10318			
2	12399	1	10318			
2	12400	1	10321			
2	12401	1	10321			
2	12402	1	10334			
2	12403	1	10334			
2	12404	1	10341			
2	12405	1	10341			
2	12406	1	10344			
2	12407	1	10344			
2	12408	1	10354			
2	12409	1	10354			
2	12410	1	10357			
2	12411	1	10357			
2	12412	1	10360			
2	12413	1	10360			
2	12414	1	10367			
2	12415	1	10367			
2	12416	1	10367			
2	12417	1	10367			
2	12418	1	10375			
2	12419	1	10375			
2	12420	1	10375			
2	12421	1	10375			
2	12422	1	10375			
2	12423	1	10381			
2	12424	1	10381			
2	12425	1	10381			
2	12426	1	10381			
2	12427	1	10381			
2	12428	1	10381			
2	12429	1	10381			
2	12430	1	10388			
2	12431	1	10388			
2	12432	1	10391			
2	12433	1	10391			
2	12434	1	10399			
2	12435	1	10399			
2	12436	1	10402			
2	12437	1	10402			
2	12438	1	10406			
2	12439	1	10406			
2	12440	1	10409			
2	12441	1	10409			
2	12442	1	10412			
2	12443	1	10412			
2	12444	1	10415			
2	12445	1	10415			
2	12446	1	10419			
2	12447	1	10419			
2	12448	1	10422			
2	12449	1	10422			
2	12450	1	10425			
2	12451	1	10425			
2	12452	1	10428			
2	12453	1	10428			
2	12454	1	2257			
2	12455	1	2257			
2	12456	1	2257			
2	12457	1	2257			
2	12458	1	2257			
2	12459	1	2257			
2	12460	1	2257			
2	12461	1	2257			
2	12462	1	2257			
2	12463	1	2257			
2	12464	1	2257			
2	12465	1	2269			
2	12466	1	2269			
2	12467	1	2269			
2	12468	1	2269			
2	12469	1	2269			
2	12470	1	2269			
2	12471	1	2287			
2	12472	1	2287			
2	12473	1	2287			
2	12474	1	2287			
2	12475	1	2287			
2	12476	1	10479			
2	12477	1	10479			
2	12478	1	10479			
2	12479	1	2293			
2	12480	1	2293			
2	12481	1	2293			
2	12482	1	2293			
2	12483	1	2293			
2	12484	1	2309			
2	12485	1	2309			
2	12486	1	2309			
2	12487	1	2309			
2	12488	1	2309			
2	12489	1	10497			
2	12490	1	10497			
2	12491	1	10497			
2	12492	1	2315			
2	12493	1	2315			
2	12494	1	2315			
2	12495	1	2315			
2	12496	1	2315			
2	12497	1	10509			
2	12498	1	10509			
2	12499	1	10512			
2	12500	1	10512			
2	12501	1	2331			
2	12502	1	2331			
2	12503	1	2331			
2	12504	1	2331			
2	12505	1	2331			
2	12506	1	10519			
2	12507	1	10519			
2	12508	1	2368			
2	12509	1	2368			
2	12510	1	2368			
2	12511	1	2368			
2	12512	1	2368			
2	12513	1	2384			
2	12514	1	2384			
2	12515	1	2384			
2	12516	1	2384			
2	12517	1	2384			
2	12518	1	2390			
2	12519	1	2390			
2	12520	1	2390			
2	12521	1	2390			
2	12522	1	2390			
2	12523	1	2406			
2	12524	1	2406			
2	12525	1	2406			
2	12526	1	2406			
2	12527	1	2406			
2	12528	1	2412			
2	12529	1	2412			
2	12530	1	2412			
2	12531	1	2412			
2	12532	1	2412			
2	12533	1	2442			
2	12534	1	2442			
2	12535	1	2442			
2	12536	1	2442			
2	12537	1	2442			
2	12538	1	2446			
2	12539	1	2446			
2	12540	1	2446			
2	12541	1	2446			
2	12542	1	2446			
2	12543	1	2450			
2	12544	1	2450			
2	12545	1	2450			
2	12546	1	2450			
2	12547	1	2450			
2	12548	1	2454			
2	12549	1	2454			
2	12550	1	2454			
2	12551	1	2454			
2	12552	1	2454			
2	12553	1	2458			
2	12554	1	2458			
2	12555	1	2458			
2	12556	1	2458			
2	12557	1	2458			
2	12558	1	2462			
2	12559	1	2462			
2	12560	1	2462			
2	12561	1	2462			
2	12562	1	2462			
2	12563	1	10652			
2	12564	1	10652			
2	12565	1	10652			
2	12566	1	10652			
2	12567	1	10652			
2	12568	1	2466			
2	12569	1	2466			
2	12570	1	2466			
2	12571	1	2466			
2	12572	1	2466			
2	12573	1	10659			
2	12574	1	10659			
2	12575	1	2470			
2	12576	1	2470			
2	12577	1	2470			
2	12578	1	2470			
2	12579	1	2470			
2	12580	1	10662			
2	12581	1	10662			
2	12582	1	10665			
2	12583	1	10665			
2	12584	1	2474			
2	12585	1	2474			
2	12586	1	2474			
2	12587	1	2474			
2	12588	1	2474			
2	12589	1	10668			
2	12590	1	10668			
2	12591	1	2478			
2	12592	1	2478			
2	12593	1	2478			
2	12594	1	2478			
2	12595	1	2478			
2	12596	1	2482			
2	12597	1	2482			
2	12598	1	2482			
2	12599	1	2482			
2	12600	1	2482			
2	12601	1	2482			
2	12602	1	2482			
2	12603	1	2482			
2	12604	1	10675			
2	12605	1	10675			
2	12606	1	10678			
2	12607	1	10678			
2	12608	1	2488			
2	12609	1	2488			
2	12610	1	2488			
2	12611	1	2488			
2	12612	1	2488			
2	12613	1	2488			
2	12614	1	2488			
2	12615	1	2488			
2	12616	1	2488			
2	12617	1	2488			
2	12618	1	2496			
2	12619	1	2496			
2	12620	1	2496			
2	12621	1	2496			
2	12622	1	2496			
2	12623	1	2496			
2	12624	1	2496			
2	12625	1	2496			
2	12626	1	10691			
2	12627	1	10691			
2	12628	1	2502			
2	12629	1	2502			
2	12630	1	2502			
2	12631	1	2502			
2	12632	1	2502			
2	12633	1	2502			
2	12634	1	2502			
2	12635	1	2502			
2	12636	1	10698			
2	12637	1	10698			
2	12638	1	2508			
2	12639	1	2508			
2	12640	1	2508			
2	12641	1	2508			
2	12642	1	2508			
2	12643	1	2508			
2	12644	1	2508			
2	12645	1	2508			
2	12646	1	10701			
2	12647	1	10701			
2	12648	1	2523			
2	12649	1	2523			
2	12650	1	2523			
2	12651	1	2523			
2	12652	1	2523			
2	12653	1	2523			
2	12654	1	2523			
2	12655	1	2533			
2	12656	1	2533			
2	12657	1	2533			
2	12658	1	2538			
2	12659	1	2538			
2	12660	1	2538			
2	12661	1	2538			
2	12662	1	2538			
2	12663	1	2542			
2	12664	1	2542			
2	12665	1	2542			
2	12666	1	2542			
2	12667	1	2542			
2	12668	1	2546			
2	12669	1	2546			
2	12670	1	2546			
2	12671	1	2546			
2	12672	1	2546			
2	12673	1	10739			
2	12674	1	10739			
2	12675	1	2550			
2	12676	1	2550			
2	12677	1	2550			
2	12678	1	2550			
2	12679	1	2550			
2	12680	1	2554			
2	12681	1	2554			
2	12682	1	2554			
2	12683	1	2554			
2	12684	1	2554			
2	12685	1	2554			
2	12686	1	2554			
2	12687	1	2554			
2	12688	1	2554			
2	12689	1	2561			
2	12690	1	2561			
2	12691	1	2561			
2	12692	1	2561			
2	12693	1	2561			
2	12694	1	2561			
2	12695	1	2561			
2	12696	1	2561			
2	12697	1	2567			
2	12698	1	2567			
2	12699	1	2567			
2	12700	1	2567			
2	12701	1	2567			
2	12702	1	2567			
2	12703	1	2567			
2	12704	1	2567			
2	12705	1	2573			
2	12706	1	2573			
2	12707	1	2573			
2	12708	1	2573			
2	12709	1	2573			
2	12710	1	2573			
2	12711	1	2573			
2	12712	1	2573			
2	12713	1	10784			
2	12714	1	10784			
2	12715	1	10784			
2	12716	1	10784			
2	12717	1	10789			
2	12718	1	10789			
2	12719	1	10792			
2	12720	1	10792			
2	12721	1	2604			
2	12722	1	2604			
2	12723	1	2604			
2	12724	1	2607			
2	12725	1	2607			
2	12726	1	2607			
2	12727	1	2607			
2	12728	1	2607			
2	12729	1	10800			
2	12730	1	10800			
2	12731	1	2611			
2	12732	1	2611			
2	12733	1	2611			
2	12734	1	2611			
2	12735	1	2611			
2	12736	1	10803			
2	12737	1	10803			
2	12738	1	10806			
2	12739	1	10806			
2	12740	1	2615			
2	12741	1	2615			
2	12742	1	2615			
2	12743	1	2615			
2	12744	1	2615			
2	12745	1	10809			
2	12746	1	10809			
2	12747	1	2619			
2	12748	1	2619			
2	12749	1	2619			
2	12750	1	2619			
2	12751	1	2619			
2	12752	1	2619			
2	12753	1	2619			
2	12754	1	2619			
2	12755	1	2619			
2	12756	1	10812			
2	12757	1	10812			
2	12758	1	10817			
2	12759	1	10817			
2	12760	1	2626			
2	12761	1	2626			
2	12762	1	2626			
2	12763	1	2626			
2	12764	1	2626			
2	12765	1	2626			
2	12766	1	2626			
2	12767	1	2626			
2	12768	1	10820			
2	12769	1	10820			
2	12770	1	2632			
2	12771	1	2632			
2	12772	1	2632			
2	12773	1	2632			
2	12774	1	2632			
2	12775	1	2632			
2	12776	1	2632			
2	12777	1	2632			
2	12778	1	2638			
2	12779	1	2638			
2	12780	1	2638			
2	12781	1	2638			
2	12782	1	2638			
2	12783	1	2638			
2	12784	1	2638			
2	12785	1	2638			
2	12786	1	2644			
2	12787	1	2644			
2	12788	1	2644			
2	12789	1	2644			
2	12790	1	2644			
2	12791	1	2644			
2	12792	1	2644			
2	12793	1	2644			
2	12794	1	2650			
2	12795	1	2650			
2	12796	1	2654			
2	12797	1	2654			
2	12798	1	2654			
2	12799	1	2654			
2	12800	1	2654			
2	12801	1	2658			
2	12802	1	2658			
2	12803	1	2658			
2	12804	1	2658			
2	12805	1	2658			
2	12806	1	2662			
2	12807	1	2662			
2	12808	1	2662			
2	12809	1	2662			
2	12810	1	2662			
2	12811	1	2666			
2	12812	1	2666			
2	12813	1	2666			
2	12814	1	2666			
2	12815	1	2666			
2	12816	1	2670			
2	12817	1	2670			
2	12818	1	2670			
2	12819	1	2670			
2	12820	1	2670			
2	12821	1	2674			
2	12822	1	2674			
2	12823	1	2674			
2	12824	1	2674			
2	12825	1	2674			
2	12826	1	2674			
2	12827	1	2674			
2	12828	1	2680			
2	12829	1	2680			
2	12830	1	2680			
2	12831	1	10876			
2	12832	1	10876			
2	12833	1	2688			
2	12834	1	2688			
2	12835	1	2688			
2	12836	1	2688			
2	12837	1	2688			
2	12838	1	10879			
2	12839	1	10879			
2	12840	1	2692			
2	12841	1	2692			
2	12842	1	2692			
2	12843	1	2692			
2	12844	1	2692			
2	12845	1	2696			
2	12846	1	2696			
2	12847	1	2696			
2	12848	1	2696			
2	12849	1	2696			
2	12850	1	2700			
2	12851	1	2700			
2	12852	1	2700			
2	12853	1	2700			
2	12854	1	2700			
2	12855	1	10892			
2	12856	1	10892			
2	12857	1	2704			
2	12858	1	2704			
2	12859	1	2704			
2	12860	1	2704			
2	12861	1	2704			
2	12862	1	10899			
2	12863	1	10899			
2	12864	1	10902			
2	12865	1	10902			
2	12866	1	2729			
2	12867	1	2729			
2	12868	1	2729			
2	12869	1	2729			
2	12870	1	2729			
2	12871	1	2733			
2	12872	1	2733			
2	12873	1	2733			
2	12874	1	2733			
2	12875	1	2733			
2	12876	1	10928			
2	12877	1	10928			
2	12878	1	2737			
2	12879	1	2737			
2	12880	1	2737			
2	12881	1	2737			
2	12882	1	2737			
2	12883	1	10931			
2	12884	1	10931			
2	12885	1	2741			
2	12886	1	2741			
2	12887	1	2741			
2	12888	1	2741			
2	12889	1	2741			
2	12890	1	2745			
2	12891	1	2745			
2	12892	1	2745			
2	12893	1	2745			
2	12894	1	2745			
2	12895	1	10938			
2	12896	1	10938			
2	12897	1	2749			
2	12898	1	2749			
2	12899	1	2749			
2	12900	1	2749			
2	12901	1	2749			
2	12902	1	10941			
2	12903	1	10941			
2	12904	1	10944			
2	12905	1	10944			
2	12906	1	2753			
2	12907	1	2753			
2	12908	1	2753			
2	12909	1	2753			
2	12910	1	2753			
2	12911	1	10947			
2	12912	1	10947			
2	12913	1	2757			
2	12914	1	2757			
2	12915	1	2757			
2	12916	1	2757			
2	12917	1	2757			
2	12918	1	10950			
2	12919	1	10950			
2	12920	1	2761			
2	12921	1	2761			
2	12922	1	2761			
2	12923	1	2761			
2	12924	1	2761			
2	12925	1	10955			
2	12926	1	10955			
2	12927	1	2766			
2	12928	1	2766			
2	12929	1	10958			
2	12930	1	10958			
2	12931	1	2769			
2	12932	1	2769			
2	12933	1	2772			
2	12934	1	2772			
2	12935	1	2775			
2	12936	1	2775			
2	12937	1	2778			
2	12938	1	2778			
2	12939	1	2781			
2	12940	1	2781			
2	12941	1	2784			
2	12942	1	2784			
2	12943	1	2787			
2	12944	1	2787			
2	12945	1	2790			
2	12946	1	2790			
2	12947	1	2793			
2	12948	1	2793			
2	12949	1	2796			
2	12950	1	2796			
2	12951	1	10992			
2	12952	1	10992			
2	12953	1	10995			
2	12954	1	10995			
2	12955	1	11008			
2	12956	1	11008			
2	12957	1	11015			
2	12958	1	11015			
2	12959	1	11018			
2	12960	1	11018			
2	12961	1	11044			
2	12962	1	11044			
2	12963	1	11047			
2	12964	1	11047			
2	12965	1	11050			
2	12966	1	11050			
2	12967	1	11053			
2	12968	1	11053			
2	12969	1	11056			
2	12970	1	11056			
2	12971	1	11059			
2	12972	1	11059			
2	12973	1	11062			
2	12974	1	11062			
2	12975	1	11067			
2	12976	1	11067			
2	12977	1	11070			
2	12978	1	11070			
2	12979	1	11100			
2	12980	1	11100			
2	12981	1	11103			
2	12982	1	11103			
2	12983	1	11124			
2	12984	1	11124			
2	12985	1	11127			
2	12986	1	11127			
2	12987	1	11130			
2	12988	1	11130			
2	12989	1	11156			
2	12990	1	11156			
2	12991	1	11159			
2	12992	1	11159			
2	12993	1	11162			
2	12994	1	11162			
2	12995	1	11165			
2	12996	1	11165			
2	12997	1	11168			
2	12998	1	11168			
2	12999	1	11171			
2	13000	1	11171			
2	13001	1	11174			
2	13002	1	11174			
2	13003	1	11177			
2	13004	1	11177			
2	13005	1	11180			
2	13006	1	11180			
2	13007	1	11205			
2	13008	1	11205			
2	13009	1	11233			
2	13010	1	11233			
2	13011	1	11236			
2	13012	1	11236			
2	13013	1	11239			
2	13014	1	11239			
2	13015	1	11252			
2	13016	1	11252			
2	13017	1	11257			
2	13018	1	11257			
2	13019	1	3073			
2	13020	1	3073			
2	13021	1	3080			
2	13022	1	3080			
2	13023	1	11272			
2	13024	1	11272			
2	13025	1	3097			
2	13026	1	3097			
2	13027	1	3097			
2	13028	1	3101			
2	13029	1	3101			
2	13030	1	3101			
2	13031	1	3101			
2	13032	1	3101			
2	13033	1	3107			
2	13034	1	3107			
2	13035	1	3107			
2	13036	1	3107			
2	13037	1	3107			
2	13038	1	3107			
2	13039	1	11299			
2	13040	1	11299			
2	13041	1	11302			
2	13042	1	11302			
2	13043	1	3114			
2	13044	1	3114			
2	13045	1	3114			
2	13046	1	3114			
2	13047	1	3114			
2	13048	1	3114			
2	13049	1	3114			
2	13050	1	3114			
2	13051	1	3122			
2	13052	1	3122			
2	13053	1	3122			
2	13054	1	3126			
2	13055	1	3126			
2	13056	1	3126			
2	13057	1	11317			
2	13058	1	11317			
2	13059	1	3131			
2	13060	1	3131			
2	13061	1	11323			
2	13062	1	11323			
2	13063	1	3137			
2	13064	1	3137			
2	13065	1	3140			
2	13066	1	3140			
2	13067	1	3140			
2	13068	1	3144			
2	13069	1	3144			
2	13070	1	3144			
2	13071	1	3144			
2	13072	1	3149			
2	13073	1	3149			
2	13074	1	3149			
2	13075	1	3149			
2	13076	1	3149			
2	13077	1	3155			
2	13078	1	3155			
2	13079	1	3155			
2	13080	1	3159			
2	13081	1	3159			
2	13082	1	3159			
2	13083	1	3169			
2	13084	1	3169			
2	13085	1	3169			
2	13086	1	3173			
2	13087	1	3173			
2	13088	1	3173			
2	13089	1	3173			
2	13090	1	3178			
2	13091	1	3178			
2	13092	1	3178			
2	13093	1	3178			
2	13094	1	3178			
2	13095	1	3178			
2	13096	1	3185			
2	13097	1	3185			
2	13098	1	3185			
2	13099	1	3189			
2	13100	1	3189			
2	13101	1	3189			
2	13102	1	3189			
2	13103	1	3189			
2	13104	1	3195			
2	13105	1	3195			
2	13106	1	3195			
2	13107	1	3195			
2	13108	1	3195			
2	13109	1	3195			
2	13110	1	3202			
2	13111	1	3202			
2	13112	1	3202			
2	13113	1	3202			
2	13114	1	3202			
2	13115	1	3202			
2	13116	1	3202			
2	13117	1	3202			
2	13118	1	3211			
2	13119	1	3211			
2	13120	1	3211			
2	13121	1	3215			
2	13122	1	3215			
2	13123	1	3215			
2	13124	1	3215			
2	13125	1	3215			
2	13126	1	3221			
2	13127	1	3221			
2	13128	1	3221			
2	13129	1	3221			
2	13130	1	3221			
2	13131	1	3221			
2	13132	1	3221			
2	13133	1	3229			
2	13134	1	3229			
2	13135	1	3232			
2	13136	1	3232			
2	13137	1	3232			
2	13138	1	3236			
2	13139	1	3236			
2	13140	1	3236			
2	13141	1	3236			
2	13142	1	3241			
2	13143	1	3241			
2	13144	1	3241			
2	13145	1	3241			
2	13146	1	3241			
2	13147	1	3247			
2	13148	1	3247			
2	13149	1	3247			
2	13150	1	3247			
2	13151	1	3247			
2	13152	1	3251			
2	13153	1	3251			
2	13154	1	3251			
2	13155	1	3251			
2	13156	1	3251			
2	13157	1	3255			
2	13158	1	3255			
2	13159	1	3255			
2	13160	1	3255			
2	13161	1	3255			
2	13162	1	3259			
2	13163	1	3259			
2	13164	1	3259			
2	13165	1	3259			
2	13166	1	3259			
2	13167	1	3263			
2	13168	1	3263			
2	13169	1	3263			
2	13170	1	3263			
2	13171	1	3263			
2	13172	1	3267			
2	13173	1	3267			
2	13174	1	3267			
2	13175	1	3267			
2	13176	1	3267			
2	13177	1	3267			
2	13178	1	3267			
2	13179	1	3267			
2	13180	1	3273			
2	13181	1	3273			
2	13182	1	3273			
2	13183	1	3273			
2	13184	1	3273			
2	13185	1	3273			
2	13186	1	3273			
2	13187	1	3273			
2	13188	1	3273			
2	13189	1	3273			
2	13190	1	3281			
2	13191	1	3281			
2	13192	1	3281			
2	13193	1	3281			
2	13194	1	3281			
2	13195	1	3281			
2	13196	1	3281			
2	13197	1	3281			
2	13198	1	3287			
2	13199	1	3287			
2	13200	1	3287			
2	13201	1	3287			
2	13202	1	3287			
2	13203	1	3287			
2	13204	1	3287			
2	13205	1	3287			
2	13206	1	3293			
2	13207	1	3293			
2	13208	1	3293			
2	13209	1	3293			
2	13210	1	3293			
2	13211	1	3293			
2	13212	1	3293			
2	13213	1	3293			
2	13214	1	3299			
2	13215	1	3299			
2	13216	1	3299			
2	13217	1	3299			
2	13218	1	3299			
2	13219	1	3303			
2	13220	1	3303			
2	13221	1	3303			
2	13222	1	3303			
2	13223	1	3303			
2	13224	1	3307			
2	13225	1	3307			
2	13226	1	3307			
2	13227	1	3307			
2	13228	1	3307			
2	13229	1	3311			
2	13230	1	3311			
2	13231	1	3311			
2	13232	1	3311			
2	13233	1	3311			
2	13234	1	3315			
2	13235	1	3315			
2	13236	1	3315			
2	13237	1	3315			
2	13238	1	3315			
2	13239	1	3315			
2	13240	1	3315			
2	13241	1	3315			
2	13242	1	3315			
2	13243	1	3322			
2	13244	1	3322			
2	13245	1	3322			
2	13246	1	3322			
2	13247	1	3322			
2	13248	1	3322			
2	13249	1	3322			
2	13250	1	3322			
2	13251	1	3328			
2	13252	1	3328			
2	13253	1	3328			
2	13254	1	3328			
2	13255	1	3328			
2	13256	1	3328			
2	13257	1	3328			
2	13258	1	3328			
2	13259	1	3334			
2	13260	1	3334			
2	13261	1	3334			
2	13262	1	3334			
2	13263	1	3334			
2	13264	1	3334			
2	13265	1	3334			
2	13266	1	3334			
2	13267	1	3340			
2	13268	1	3340			
2	13269	1	3340			
2	13270	1	3343			
2	13271	1	3343			
2	13272	1	3343			
2	13273	1	3343			
2	13274	1	3343			
2	13275	1	3343			
2	13276	1	3343			
2	13277	1	3343			
2	13278	1	3349			
2	13279	1	3349			
2	13280	1	3349			
2	13281	1	3349			
2	13282	1	3349			
2	13283	1	3349			
2	13284	1	3349			
2	13285	1	3349			
2	13286	1	3355			
2	13287	1	3355			
2	13288	1	3355			
2	13289	1	3355			
2	13290	1	3355			
2	13291	1	3355			
2	13292	1	3355			
2	13293	1	3355			
2	13294	1	3375			
2	13295	1	3375			
2	13296	1	3375			
2	13297	1	3381			
2	13298	1	3381			
2	13299	1	3381			
2	13300	1	3384			
2	13301	1	3384			
2	13302	1	3384			
2	13303	1	3384			
2	13304	1	3384			
2	13305	1	3384			
2	13306	1	3384			
2	13307	1	3384			
2	13308	1	3390			
2	13309	1	3390			
2	13310	1	3390			
2	13311	1	3390			
2	13312	1	3390			
2	13313	1	3390			
2	13314	1	3390			
2	13315	1	3390			
2	13316	1	3390			
2	13317	1	3390			
2	13318	1	3398			
2	13319	1	3398			
2	13320	1	3398			
2	13321	1	3398			
2	13322	1	3398			
2	13323	1	3398			
2	13324	1	3398			
2	13325	1	3398			
2	13326	1	3404			
2	13327	1	3404			
2	13328	1	3404			
2	13329	1	3404			
2	13330	1	3404			
2	13331	1	3404			
2	13332	1	3404			
2	13333	1	3404			
2	13334	1	3410			
2	13335	1	3410			
2	13336	1	3410			
2	13337	1	3410			
2	13338	1	3410			
2	13339	1	3410			
2	13340	1	3410			
2	13341	1	3410			
2	13342	1	3416			
2	13343	1	3416			
2	13344	1	3416			
2	13345	1	3416			
2	13346	1	3416			
2	13347	1	3420			
2	13348	1	3420			
2	13349	1	3420			
2	13350	1	3420			
2	13351	1	3420			
2	13352	1	3424			
2	13353	1	3424			
2	13354	1	3424			
2	13355	1	3424			
2	13356	1	3424			
2	13357	1	3428			
2	13358	1	3428			
2	13359	1	3428			
2	13360	1	3428			
2	13361	1	3428			
2	13362	1	3432			
2	13363	1	3432			
2	13364	1	3432			
2	13365	1	3432			
2	13366	1	3432			
2	13367	1	3436			
2	13368	1	3436			
2	13369	1	3436			
2	13370	1	3436			
2	13371	1	3436			
2	13372	1	3440			
2	13373	1	3440			
2	13374	1	3440			
2	13375	1	3440			
2	13376	1	3440			
2	13377	1	3444			
2	13378	1	3444			
2	13379	1	3444			
2	13380	1	3444			
2	13381	1	3444			
2	13382	1	3448			
2	13383	1	3448			
2	13384	1	3448			
2	13385	1	3448			
2	13386	1	3448			
2	13387	1	3454			
2	13388	1	3454			
2	13389	1	3454			
2	13390	1	3454			
2	13391	1	3454			
2	13392	1	3458			
2	13393	1	3458			
2	13394	1	3458			
2	13395	1	3458			
2	13396	1	3458			
2	13397	1	3462			
2	13398	1	3462			
2	13399	1	3462			
2	13400	1	3462			
2	13401	1	3462			
2	13402	1	3466			
2	13403	1	3466			
2	13404	1	3466			
2	13405	1	3466			
2	13406	1	3466			
2	13407	1	3470			
2	13408	1	3470			
2	13409	1	3470			
2	13410	1	3470			
2	13411	1	3470			
2	13412	1	3474			
2	13413	1	3474			
2	13414	1	3474			
2	13415	1	3474			
2	13416	1	3474			
2	13417	1	3478			
2	13418	1	3478			
2	13419	1	3478			
2	13420	1	3478			
2	13421	1	3478			
2	13422	1	3482			
2	13423	1	3482			
2	13424	1	3482			
2	13425	1	3482			
2	13426	1	3482			
2	13427	1	3507			
2	13428	1	3507			
2	13429	1	3515			
2	13430	1	3515			
2	13431	1	3625			
2	13432	1	3625			
2	13433	1	3628			
2	13434	1	3628			
2	13435	1	3658			
2	13436	1	3658			
2	13437	1	3783			
2	13438	1	3783			
2	13439	1	3786			
2	13440	1	3786			
2	13441	1	10522			
2	13442	1	10522			
2	13443	1	3789			
2	13444	1	3789			
2	13445	1	10525			
2	13446	1	10525			
2	13447	1	10528			
2	13448	1	10528			
2	13449	1	10531			
2	13450	1	10531			
2	13451	1	10536			
2	13452	1	10536			
2	13453	1	10539			
2	13454	1	10539			
2	13455	1	3885			
2	13456	1	3885			
2	13457	1	3888			
2	13458	1	3888			
2	13459	1	3891			
2	13460	1	3891			
2	13461	1	10583			
2	13462	1	10583			
2	13463	1	10583			
2	13464	1	10589			
2	13465	1	10589			
2	13466	1	10589			
2	13467	1	10589			
2	13468	1	4193			
2	13469	1	4193			
2	13470	1	4193			
2	13471	1	4303			
2	13472	1	4303			
2	13473	1	4545			
2	13474	1	4545			
2	13475	1	4545			
2	13476	1	4549			
2	13477	1	4549			
2	13478	1	4549			
2	13479	1	4549			
2	13480	1	4549			
2	13481	1	4555			
2	13482	1	4555			
2	13483	1	4555			
2	13484	1	4555			
2	13485	1	4555			
2	13486	1	4555			
2	13487	1	4555			
2	13488	1	4563			
2	13489	1	4563			
2	13490	1	4566			
2	13491	1	4566			
2	13492	1	4566			
2	13493	1	4570			
2	13494	1	4570			
2	13495	1	4570			
2	13496	1	4570			
2	13497	1	4577			
2	13498	1	4577			
2	13499	1	4577			
2	13500	1	4581			
2	13501	1	4581			
2	13502	1	4581			
2	13503	1	4581			
2	13504	1	4586			
2	13505	1	4586			
2	13506	1	4586			
2	13507	1	4586			
2	13508	1	4586			
2	13509	1	4586			
2	13510	1	4593			
2	13511	1	4593			
2	13512	1	4593			
2	13513	1	4597			
2	13514	1	4597			
2	13515	1	4597			
2	13516	1	4597			
2	13517	1	4597			
2	13518	1	4603			
2	13519	1	4603			
2	13520	1	4603			
2	13521	1	4603			
2	13522	1	4603			
2	13523	1	4603			
2	13524	1	4657			
2	13525	1	4657			
2	13526	1	4657			
2	13527	1	4661			
2	13528	1	4661			
2	13529	1	4661			
2	13530	1	4661			
2	13531	1	4661			
2	13532	1	4667			
2	13533	1	4667			
2	13534	1	4667			
2	13535	1	4667			
2	13536	1	4667			
2	13537	1	4667			
2	13538	1	4667			
2	13539	1	4675			
2	13540	1	4675			
2	13541	1	4678			
2	13542	1	4678			
2	13543	1	4678			
2	13544	1	4682			
2	13545	1	4682			
2	13546	1	4682			
2	13547	1	4682			
2	13548	1	4687			
2	13549	1	4687			
2	13550	1	4687			
2	13551	1	4687			
2	13552	1	4687			
2	13553	1	4702			
2	13554	1	4702			
2	13555	1	4702			
2	13556	1	4706			
2	13557	1	4706			
2	13558	1	4706			
2	13559	1	4706			
2	13560	1	4711			
2	13561	1	4711			
2	13562	1	4711			
2	13563	1	4711			
2	13564	1	4711			
2	13565	1	4711			
2	13566	1	4718			
2	13567	1	4718			
2	13568	1	4718			
2	13569	1	4722			
2	13570	1	4722			
2	13571	1	4722			
2	13572	1	4722			
2	13573	1	4722			
2	13574	1	4728			
2	13575	1	4728			
2	13576	1	4728			
2	13577	1	4728			
2	13578	1	4728			
2	13579	1	4728			
2	13580	1	4735			
2	13581	1	4735			
2	13582	1	4735			
2	13583	1	4735			
2	13584	1	4735			
2	13585	1	4735			
2	13586	1	4735			
2	13587	1	4735			
2	13588	1	4769			
2	13589	1	4769			
2	13590	1	4769			
2	13591	1	4769			
2	13592	1	4769			
2	13593	1	4769			
2	13594	1	4769			
2	13595	1	4784			
2	13596	1	4784			
2	13597	1	4790			
2	13598	1	4790			
2	13599	1	4803			
2	13600	1	4803			
2	13601	1	4806			
2	13602	1	4806			
2	13603	1	4844			
2	13604	1	4844			
2	13605	1	4871			
2	13606	1	4871			
2	13607	1	4940			
2	13608	1	4940			
2	13609	1	4997			
2	13610	1	4997			
2	13611	1	5027			
2	13612	1	5027			
2	13613	1	5030			
2	13614	1	5030			
2	13615	1	5632			
2	13616	1	5632			
2	13617	1	5632			
2	13618	1	5632			
2	13619	1	5632			
2	13620	1	5632			
2	13621	1	5632			
2	13622	1	5632			
2	13623	1	5632			
2	13624	1	5640			
2	13625	1	5640			
2	13626	1	5640			
2	13627	1	5640			
2	13628	1	5640			
2	13629	1	5640			
2	13630	1	5640			
2	13631	1	5640			
2	13632	1	5640			
2	13633	1	5640			
2	13634	1	5640			
2	13635	1	5640			
2	13636	1	5640			
2	13637	1	5640			
2	13638	1	5640			
2	13639	1	5654			
2	13640	1	5654			
2	13641	1	5654			
2	13642	1	5654			
2	13643	1	5654			
2	13644	1	5654			
2	13645	1	5654			
2	13646	1	5654			
2	13647	1	5654			
2	13648	1	5654			
2	13649	1	5654			
2	13650	1	5654			
2	13651	1	5654			
2	13652	1	5654			
2	13653	1	5654			
2	13654	1	5654			
2	13655	1	5654			
2	13656	1	5670			
2	13657	1	5670			
2	13658	1	5670			
2	13659	1	5670			
2	13660	1	5670			
2	13661	1	5670			
2	13662	1	5670			
2	13663	1	5670			
2	13664	1	5670			
2	13665	1	5670			
2	13666	1	5670			
2	13667	1	5670			
2	13668	1	5670			
2	13669	1	5670			
2	13670	1	5683			
2	13671	1	5683			
2	13672	1	5683			
2	13673	1	5683			
2	13674	1	5683			
2	13675	1	5683			
2	13676	1	5683			
2	13677	1	5683			
2	13678	1	5690			
2	13679	1	5690			
2	13680	1	5690			
2	13681	1	5690			
2	13682	1	5690			
2	13683	1	5690			
2	13684	1	5690			
2	13685	1	5697			
2	13686	1	5697			
2	13687	1	5697			
2	13688	1	5697			
2	13689	1	5697			
2	13690	1	5697			
2	13691	1	5697			
2	13692	1	5697			
2	13693	1	5697			
2	13694	1	5697			
2	13695	1	5707			
2	13696	1	5707			
2	13697	1	5707			
2	13698	1	5707			
2	13699	1	5707			
2	13700	1	5707			
2	13701	1	5707			
2	13702	1	5707			
2	13703	1	5707			
2	13704	1	5707			
2	13705	1	5707			
2	13706	1	5718			
2	13707	1	5718			
2	13708	1	5718			
2	13709	1	5718			
2	13710	1	5718			
2	13711	1	5718			
2	13712	1	5718			
2	13713	1	5718			
2	13714	1	5718			
2	13715	1	5718			
2	13716	1	5728			
2	13717	1	5728			
2	13718	1	5728			
2	13719	1	5728			
2	13720	1	5728			
2	13721	1	5728			
2	13722	1	5728			
2	13723	1	5736			
2	13724	1	5736			
2	13725	1	5736			
2	13726	1	5740			
2	13727	1	5740			
2	13728	1	5740			
2	13729	1	5744			
2	13730	1	5744			
2	13731	1	5744			
2	13732	1	5744			
2	13733	1	5747			
2	13734	1	5747			
2	13735	1	5747			
2	13736	1	5751			
2	13737	1	5751			
2	13738	1	5751			
2	13739	1	5755			
2	13740	1	5755			
2	13741	1	5755			
2	13742	1	5755			
2	13743	1	5758			
2	13744	1	5758			
2	13745	1	5758			
2	13746	1	5762			
2	13747	1	5762			
2	13748	1	5762			
2	13749	1	5766			
2	13750	1	5766			
2	13751	1	5766			
2	13752	1	5766			
2	13753	1	5771			
2	13754	1	5771			
2	13755	1	5771			
2	13756	1	5771			
2	13757	1	5771			
2	13758	1	5771			
2	13759	1	5771			
2	13760	1	5771			
2	13761	1	5778			
2	13762	1	5778			
2	13763	1	5778			
2	13764	1	5778			
2	13765	1	5778			
2	13766	1	5778			
2	13767	1	5778			
2	13768	1	5778			
2	13769	1	5778			
2	13770	1	5778			
2	13771	1	5778			
2	13772	1	5778			
2	13773	1	5789			
2	13774	1	5789			
2	13775	1	5789			
2	13776	1	5789			
2	13777	1	5789			
2	13778	1	5789			
2	13779	1	5789			
2	13780	1	5789			
2	13781	1	5789			
2	13782	1	5789			
2	13783	1	5789			
2	13784	1	5799			
2	13785	1	5799			
2	13786	1	5799			
2	13787	1	5799			
2	13788	1	5799			
2	13789	1	5799			
2	13790	1	5799			
2	13791	1	5799			
2	13792	1	5799			
2	13793	1	5807			
2	13794	1	5807			
2	13795	1	5807			
2	13796	1	5807			
2	13797	1	5807			
2	13798	1	5807			
2	13799	1	5807			
2	13800	1	5807			
2	13801	1	5807			
2	13802	1	5807			
2	13803	1	5807			
2	13804	1	5807			
2	13805	1	5807			
2	13806	1	5807			
2	13807	1	5807			
2	13808	1	5821			
2	13809	1	5821			
2	13810	1	5821			
2	13811	1	5821			
2	13812	1	5821			
2	13813	1	5821			
2	13814	1	5821			
2	13815	1	5821			
2	13816	1	5821			
2	13817	1	5821			
2	13818	1	5821			
2	13819	1	5821			
2	13820	1	5821			
2	13821	1	5821			
2	13822	1	5821			
2	13823	1	5821			
2	13824	1	5821			
2	13825	1	5837			
2	13826	1	5837			
2	13827	1	5837			
2	13828	1	5837			
2	13829	1	5837			
2	13830	1	5837			
2	13831	1	5837			
2	13832	1	5837			
2	13833	1	5837			
2	13834	1	5837			
2	13835	1	5837			
2	13836	1	5837			
2	13837	1	5837			
2	13838	1	5837			
2	13839	1	10141			
2	13840	1	10141			
2	13841	1	10141			
2	13842	1	10141			
2	13843	1	10141			
2	13844	1	10141			
2	13845	1	10141			
2	13846	1	5850			
2	13847	1	5850			
2	13848	1	5850			
2	13849	1	5850			
2	13850	1	5850			
2	13851	1	5850			
2	13852	1	5850			
2	13853	1	5856			
2	13854	1	5856			
2	13855	1	5856			
2	13856	1	5856			
2	13857	1	5856			
2	13858	1	5856			
2	13859	1	5856			
2	13860	1	5856			
2	13861	1	5863			
2	13862	1	5863			
2	13863	1	5863			
2	13864	1	5863			
2	13865	1	5863			
2	13866	1	5863			
2	13867	1	5863			
2	13868	1	5863			
2	13869	1	5870			
2	13870	1	5870			
2	13871	1	5870			
2	13872	1	5870			
2	13873	1	5870			
2	13874	1	5870			
2	13875	1	5870			
2	13876	1	5870			
2	13877	1	5870			
2	13878	1	5870			
2	13879	1	5870			
2	13880	1	5870			
2	13881	1	5881			
2	13882	1	5881			
2	13883	1	5881			
2	13884	1	5881			
2	13885	1	5881			
2	13886	1	5881			
2	13887	1	5881			
2	13888	1	5881			
2	13889	1	5881			
2	13890	1	5881			
2	13891	1	5881			
2	13892	1	5881			
2	13893	1	10003			
2	13894	1	10003			
2	13895	1	5892			
2	13896	1	5892			
2	13897	1	5892			
2	13898	1	5892			
2	13899	1	5892			
2	13900	1	5898			
2	13901	1	5898			
2	13902	1	5898			
2	13903	1	5898			
2	13904	1	5898			
2	13905	1	5898			
2	13906	1	5898			
2	13907	1	5905			
2	13908	1	5905			
2	13909	1	5905			
2	13910	1	5905			
2	13911	1	5905			
2	13912	1	5905			
2	13913	1	5905			
2	13914	1	5905			
2	13915	1	5905			
2	13916	1	5905			
2	13917	1	5915			
2	13918	1	5915			
2	13919	1	5915			
2	13920	1	5915			
2	13921	1	5915			
2	13922	1	5915			
2	13923	1	5915			
2	13924	1	5915			
2	13925	1	5915			
2	13926	1	5915			
2	13927	1	5915			
2	13928	1	5926			
2	13929	1	5926			
2	13930	1	5926			
2	13931	1	5926			
2	13932	1	5926			
2	13933	1	5926			
2	13934	1	5926			
2	13935	1	5926			
2	13936	1	5926			
2	13937	1	5926			
2	13938	1	5936			
2	13939	1	5936			
2	13940	1	5936			
2	13941	1	5936			
2	13942	1	5936			
2	13943	1	5936			
2	13944	1	5936			
2	13945	1	5960			
2	13946	1	5960			
2	13947	1	5960			
2	13948	1	5960			
2	13949	1	5960			
2	13950	1	5981			
2	13951	1	5981			
2	13952	1	5981			
2	13953	1	5981			
2	13954	1	5981			
2	13955	1	5981			
2	13956	1	5981			
2	13957	1	5981			
2	13958	1	5991			
2	13959	1	5991			
2	13960	1	5991			
2	13961	1	5991			
2	13962	1	5996			
2	13963	1	5996			
2	13964	1	5996			
2	13965	1	6000			
2	13966	1	6000			
2	13967	1	6003			
2	13968	1	6003			
2	13969	1	6003			
2	13970	1	6003			
2	13971	1	6003			
2	13972	1	6009			
2	13973	1	6009			
2	13974	1	6009			
2	13975	1	6009			
2	13976	1	6014			
2	13977	1	6014			
2	13978	1	6014			
2	13979	1	6018			
2	13980	1	6018			
2	13981	1	6041			
2	13982	1	6041			
2	13983	1	6041			
2	13984	1	6041			
2	13985	1	6041			
2	13986	1	6047			
2	13987	1	6047			
2	13988	1	6047			
2	13989	1	6047			
2	13990	1	6052			
2	13991	1	6052			
2	13992	1	6052			
2	13993	1	6056			
2	13994	1	6056			
2	13995	1	6079			
2	13996	1	6079			
2	13997	1	6079			
2	13998	1	6083			
2	13999	1	6083			
2	14000	1	6083			
2	14001	1	6087			
2	14002	1	6087			
2	14003	1	6087			
2	14004	1	6087			
2	14005	1	6127			
2	14006	1	6127			
2	14007	1	6127			
2	14008	1	6131			
2	14009	1	6131			
2	14010	1	6131			
2	14011	1	6137			
2	14012	1	6137			
2	14013	1	6137			
2	14014	1	6141			
2	14015	1	6141			
2	14016	1	6141			
2	14017	1	6145			
2	14018	1	6145			
2	14019	1	6145			
2	14020	1	6145			
2	14021	1	6166			
2	14022	1	6166			
2	14023	1	6166			
2	14024	1	6170			
2	14025	1	6170			
2	14026	1	6170			
2	14027	1	6174			
2	14028	1	6174			
2	14029	1	6174			
2	14030	1	6174			
2	14031	1	6177			
2	14032	1	6177			
2	14033	1	6177			
2	14034	1	6196			
2	14035	1	6196			
2	14036	1	6199			
2	14037	1	6199			
2	14038	1	6217			
2	14039	1	6217			
2	14040	1	6243			
2	14041	1	6243			
2	14042	1	6246			
2	14043	1	6246			
2	14044	1	6249			
2	14045	1	6249			
2	14046	1	6252			
2	14047	1	6252			
2	14048	1	6263			
2	14049	1	6263			
2	14050	1	6266			
2	14051	1	6266			
2	14052	1	6762			
2	14053	1	6762			
2	14054	1	6762			
2	14055	1	6784			
2	14056	1	6784			
2	14057	1	6797			
2	14058	1	6797			
2	14059	1	6800			
2	14060	1	6800			
2	14061	1	6803			
2	14062	1	6803			
2	14063	1	6806			
2	14064	1	6806			
2	14065	1	6809			
2	14066	1	6809			
2	14067	1	6812			
2	14068	1	6812			
2	14069	1	6833			
2	14070	1	6833			
2	14071	1	6845			
2	14072	1	6845			
2	14073	1	6867			
2	14074	1	6867			
2	14075	1	6881			
2	14076	1	6881			
2	14077	1	6894			
2	14078	1	6894			
2	14079	1	6894			
2	14080	1	6894			
2	14081	1	6894			
2	14082	1	6894			
2	14083	1	6894			
2	14084	1	6894			
2	14085	1	6901			
2	14086	1	6901			
2	14087	1	6901			
2	14088	1	6901			
2	14089	1	6901			
2	14090	1	6901			
2	14091	1	6901			
2	14092	1	6901			
2	14093	1	6901			
2	14094	1	6901			
2	14095	1	6901			
2	14096	1	6901			
2	14097	1	6912			
2	14098	1	6912			
2	14099	1	6912			
2	14100	1	6912			
2	14101	1	6912			
2	14102	1	6912			
2	14103	1	6912			
2	14104	1	6912			
2	14105	1	6912			
2	14106	1	6912			
2	14107	1	6912			
2	14108	1	6912			
2	14109	1	6923			
2	14110	1	6923			
2	14111	1	6923			
2	14112	1	6923			
2	14113	1	6923			
2	14114	1	6929			
2	14115	1	6929			
2	14116	1	6929			
2	14117	1	6929			
2	14118	1	6929			
2	14119	1	6929			
2	14120	1	6929			
2	14121	1	6936			
2	14122	1	6936			
2	14123	1	6936			
2	14124	1	6936			
2	14125	1	6936			
2	14126	1	6936			
2	14127	1	6936			
2	14128	1	6936			
2	14129	1	6936			
2	14130	1	6936			
2	14131	1	6946			
2	14132	1	6946			
2	14133	1	6946			
2	14134	1	6946			
2	14135	1	6946			
2	14136	1	6946			
2	14137	1	6946			
2	14138	1	6946			
2	14139	1	6946			
2	14140	1	6946			
2	14141	1	6946			
2	14142	1	6957			
2	14143	1	6957			
2	14144	1	6957			
2	14145	1	6957			
2	14146	1	6957			
2	14147	1	6957			
2	14148	1	6957			
2	14149	1	6957			
2	14150	1	6957			
2	14151	1	6957			
2	14152	1	6970			
2	14153	1	6970			
2	14154	1	6970			
2	14155	1	6970			
2	14156	1	6970			
2	14157	1	6970			
2	14158	1	6970			
2	14159	1	6970			
2	14160	1	6977			
2	14161	1	6977			
2	14162	1	6977			
2	14163	1	6977			
2	14164	1	6977			
2	14165	1	6977			
2	14166	1	6977			
2	14167	1	6977			
2	14168	1	6977			
2	14169	1	6977			
2	14170	1	6977			
2	14171	1	6977			
2	14172	1	6988			
2	14173	1	6988			
2	14174	1	6988			
2	14175	1	6988			
2	14176	1	6988			
2	14177	1	6988			
2	14178	1	6988			
2	14179	1	6988			
2	14180	1	6988			
2	14181	1	6988			
2	14182	1	6988			
2	14183	1	6998			
2	14184	1	6998			
2	14185	1	6998			
2	14186	1	6998			
2	14187	1	6998			
2	14188	1	6998			
2	14189	1	6998			
2	14190	1	6998			
2	14191	1	6998			
2	14192	1	7006			
2	14193	1	7006			
2	14194	1	7006			
2	14195	1	7006			
2	14196	1	7006			
2	14197	1	7006			
2	14198	1	7006			
2	14199	1	7006			
2	14200	1	7006			
2	14201	1	7006			
2	14202	1	7006			
2	14203	1	7006			
2	14204	1	7006			
2	14205	1	7006			
2	14206	1	7006			
2	14207	1	7020			
2	14208	1	7020			
2	14209	1	7020			
2	14210	1	7020			
2	14211	1	7020			
2	14212	1	7020			
2	14213	1	7020			
2	14214	1	7020			
2	14215	1	7020			
2	14216	1	7020			
2	14217	1	7020			
2	14218	1	7020			
2	14219	1	7020			
2	14220	1	7020			
2	14221	1	7020			
2	14222	1	7020			
2	14223	1	7020			
2	14224	1	7036			
2	14225	1	7036			
2	14226	1	7036			
2	14227	1	7036			
2	14228	1	7036			
2	14229	1	7036			
2	14230	1	7036			
2	14231	1	7036			
2	14232	1	7036			
2	14233	1	7036			
2	14234	1	7036			
2	14235	1	7036			
2	14236	1	7036			
2	14237	1	7036			
2	14238	1	7049			
2	14239	1	7049			
2	14240	1	7049			
2	14241	1	7049			
2	14242	1	7049			
2	14243	1	7049			
2	14244	1	7049			
2	14245	1	7057			
2	14246	1	7057			
2	14247	1	7068			
2	14248	1	7068			
2	14249	1	7068			
2	14250	1	7068			
2	14251	1	7073			
2	14252	1	7073			
2	14253	1	7073			
2	14254	1	7077			
2	14255	1	7077			
2	14256	1	7080			
2	14257	1	7080			
2	14258	1	7080			
2	14259	1	7080			
2	14260	1	7080			
2	14261	1	7086			
2	14262	1	7086			
2	14263	1	7086			
2	14264	1	7086			
2	14265	1	7091			
2	14266	1	7091			
2	14267	1	7091			
2	14268	1	7095			
2	14269	1	7095			
2	14270	1	7100			
2	14271	1	7100			
2	14272	1	7107			
2	14273	1	7107			
2	14274	1	7107			
2	14275	1	7107			
2	14276	1	7107			
2	14277	1	7107			
2	14278	1	7107			
2	14279	1	7107			
2	14280	1	7114			
2	14281	1	7114			
2	14282	1	7114			
2	14283	1	7114			
2	14284	1	7114			
2	14285	1	7114			
2	14286	1	7114			
2	14287	1	7114			
2	14288	1	7114			
2	14289	1	7114			
2	14290	1	7114			
2	14291	1	7114			
2	14292	1	7125			
2	14293	1	7125			
2	14294	1	7125			
2	14295	1	7125			
2	14296	1	7125			
2	14297	1	7125			
2	14298	1	7125			
2	14299	1	7125			
2	14300	1	7125			
2	14301	1	7125			
2	14302	1	7125			
2	14303	1	7125			
2	14304	1	7136			
2	14305	1	7136			
2	14306	1	7136			
2	14307	1	7136			
2	14308	1	7136			
2	14309	1	7142			
2	14310	1	7142			
2	14311	1	7142			
2	14312	1	7142			
2	14313	1	7142			
2	14314	1	7142			
2	14315	1	7142			
2	14316	1	7149			
2	14317	1	7149			
2	14318	1	7149			
2	14319	1	7149			
2	14320	1	7149			
2	14321	1	7149			
2	14322	1	7149			
2	14323	1	7149			
2	14324	1	7149			
2	14325	1	7149			
2	14326	1	7159			
2	14327	1	7159			
2	14328	1	7159			
2	14329	1	7159			
2	14330	1	7159			
2	14331	1	7159			
2	14332	1	7159			
2	14333	1	7159			
2	14334	1	7159			
2	14335	1	7159			
2	14336	1	7159			
2	14337	1	7170			
2	14338	1	7170			
2	14339	1	7170			
2	14340	1	7170			
2	14341	1	7170			
2	14342	1	7170			
2	14343	1	7170			
2	14344	1	7170			
2	14345	1	7170			
2	14346	1	7170			
2	14347	1	7180			
2	14348	1	7180			
2	14349	1	7180			
2	14350	1	7180			
2	14351	1	7180			
2	14352	1	7180			
2	14353	1	7180			
2	14354	1	7188			
2	14355	1	7188			
2	14356	1	7191			
2	14357	1	7191			
2	14358	1	7194			
2	14359	1	7194			
2	14360	1	7194			
2	14361	1	7198			
2	14362	1	7198			
2	14363	1	7198			
2	14364	1	7202			
2	14365	1	7202			
2	14366	1	7202			
2	14367	1	7202			
2	14368	1	7205			
2	14369	1	7205			
2	14370	1	7205			
2	14371	1	7209			
2	14372	1	7209			
2	14373	1	7209			
2	14374	1	7213			
2	14375	1	7213			
2	14376	1	7213			
2	14377	1	7213			
2	14378	1	7222			
2	14379	1	7222			
2	14380	1	7222			
2	14381	1	7222			
2	14382	1	7222			
2	14383	1	7222			
2	14384	1	7222			
2	14385	1	7222			
2	14386	1	7229			
2	14387	1	7229			
2	14388	1	7229			
2	14389	1	7229			
2	14390	1	7229			
2	14391	1	7229			
2	14392	1	7229			
2	14393	1	7229			
2	14394	1	7229			
2	14395	1	7229			
2	14396	1	7229			
2	14397	1	7229			
2	14398	1	7240			
2	14399	1	7240			
2	14400	1	7240			
2	14401	1	7240			
2	14402	1	7240			
2	14403	1	7240			
2	14404	1	7240			
2	14405	1	7240			
2	14406	1	7240			
2	14407	1	7240			
2	14408	1	7240			
2	14409	1	7250			
2	14410	1	7250			
2	14411	1	7250			
2	14412	1	7250			
2	14413	1	7250			
2	14414	1	7250			
2	14415	1	7250			
2	14416	1	7250			
2	14417	1	7250			
2	14418	1	7258			
2	14419	1	7258			
2	14420	1	7258			
2	14421	1	7258			
2	14422	1	7258			
2	14423	1	7258			
2	14424	1	7258			
2	14425	1	7258			
2	14426	1	7258			
2	14427	1	7258			
2	14428	1	7258			
2	14429	1	7258			
2	14430	1	7258			
2	14431	1	7258			
2	14432	1	7258			
2	14433	1	7272			
2	14434	1	7272			
2	14435	1	7272			
2	14436	1	7272			
2	14437	1	7272			
2	14438	1	7272			
2	14439	1	7272			
2	14440	1	7272			
2	14441	1	7272			
2	14442	1	7272			
2	14443	1	7272			
2	14444	1	7272			
2	14445	1	7272			
2	14446	1	7272			
2	14447	1	7272			
2	14448	1	7272			
2	14449	1	7272			
2	14450	1	7288			
2	14451	1	7288			
2	14452	1	7288			
2	14453	1	7288			
2	14454	1	7288			
2	14455	1	7288			
2	14456	1	7288			
2	14457	1	7288			
2	14458	1	7288			
2	14459	1	7288			
2	14460	1	7288			
2	14461	1	7288			
2	14462	1	7288			
2	14463	1	7288			
2	14464	1	7301			
2	14465	1	7301			
2	14466	1	7301			
2	14467	1	7301			
2	14468	1	7301			
2	14469	1	7301			
2	14470	1	7301			
2	14471	1	7307			
2	14472	1	7307			
2	14473	1	7307			
2	14474	1	7307			
2	14475	1	7307			
2	14476	1	7307			
2	14477	1	7307			
2	14478	1	7307			
2	14479	1	7314			
2	14480	1	7314			
2	14481	1	7314			
2	14482	1	7318			
2	14483	1	7318			
2	14484	1	7318			
2	14485	1	7322			
2	14486	1	7322			
2	14487	1	7322			
2	14488	1	7322			
2	14489	1	7325			
2	14490	1	7325			
2	14491	1	7328			
2	14492	1	7328			
2	14493	1	7331			
2	14494	1	7331			
2	14495	1	7331			
2	14496	1	7331			
2	14497	1	7334			
2	14498	1	7334			
2	14499	1	7337			
2	14500	1	7337			
2	14501	1	7346			
2	14502	1	7346			
2	14503	1	7346			
2	14504	1	7346			
2	14505	1	7351			
2	14506	1	7351			
2	14507	1	7351			
2	14508	1	7355			
2	14509	1	7355			
2	14510	1	7358			
2	14511	1	7358			
2	14512	1	7358			
2	14513	1	7358			
2	14514	1	7358			
2	14515	1	7364			
2	14516	1	7364			
2	14517	1	7364			
2	14518	1	7364			
2	14519	1	7369			
2	14520	1	7369			
2	14521	1	7369			
2	14522	1	7373			
2	14523	1	7373			
2	14524	1	7378			
2	14525	1	7378			
2	14526	1	7381			
2	14527	1	7381			
2	14528	1	7384			
2	14529	1	7384			
2	14530	1	7387			
2	14531	1	7387			
2	14532	1	7387			
2	14533	1	7391			
2	14534	1	7391			
2	14535	1	7391			
2	14536	1	7391			
2	14537	1	7394			
2	14538	1	7394			
2	14539	1	7394			
2	14540	1	7398			
2	14541	1	7398			
2	14542	1	7398			
2	14543	1	7402			
2	14544	1	7402			
2	14545	1	7402			
2	14546	1	7402			
2	14547	1	7441			
2	14548	1	7441			
2	14549	1	7444			
2	14550	1	7444			
2	14551	1	7560			
2	14552	1	7560			
2	14553	1	7563			
2	14554	1	7563			
2	14555	1	7566			
2	14556	1	7566			
2	14557	1	7569			
2	14558	1	7569			
2	14559	1	7574			
2	14560	1	7574			
2	14561	1	7577			
2	14562	1	7577			
2	14563	1	7582			
2	14564	1	7582			
2	14565	1	7585			
2	14566	1	7585			
2	14567	1	7588			
2	14568	1	7588			
2	14569	1	7591			
2	14570	1	7591			
2	14571	1	7609			
2	14572	1	7609			
2	14573	1	7609			
2	14574	1	7613			
2	14575	1	7613			
2	14576	1	7620			
2	14577	1	7620			
2	14578	1	7650			
2	14579	1	7650			
2	14580	1	7655			
2	14581	1	7655			
2	14582	1	7655			
2	14583	1	7659			
2	14584	1	7659			
2	14585	1	7671			
2	14586	1	7671			
2	14587	1	7852			
2	14588	1	7852			
2	14589	1	8114			
2	14590	1	8114			
2	14591	1	8117			
2	14592	1	8117			
2	14593	1	8131			
2	14594	1	8131			
2	14595	1	8134			
2	14596	1	8134			
2	14597	1	8146			
2	14598	1	8146			
2	14599	1	8156			
2	14600	1	8156			
2	14601	1	8166			
2	14602	1	8166			
2	14603	1	8169			
2	14604	1	8169			
2	14605	1	8183			
2	14606	1	8183			
2	14607	1	8186			
2	14608	1	8186			
