1 1 0 6 0
1 8 0 4 0
1 13 0 3 0
1 17 0 8 0
1 26 0 2 0
1 29 0 6 0
1 36 0 5 0
1 42 0 8 0
1 51 0 3 0
1 55 0 3 0
1 59 0 8 0
1 68 0 3 0
1 72 0 1 0
1 73 0 1 0
1 74 0 1 0
1 75 0 4 0
1 80 0 4 0
1 85 0 1 0
1 86 0 1 0
1 87 0 1 0
1 88 0 1 0
1 89 0 1 0
1 90 0 1 0
1 91 0 4 0
1 96 0 4 0
1 101 0 4 0
1 106 0 4 0
1 111 0 4 0
1 116 0 4 0
1 121 0 4 0
1 126 0 3 0
1 130 0 4 0
1 135 0 2 0
1 138 0 4 0
1 143 0 2 0
1 146 0 2 0
1 149 0 2 0
1 152 0 1 0
1 153 0 2 0
1 156 0 2 0
1 159 0 5 0
1 165 0 5 0
1 171 0 5 0
1 177 0 5 0
1 183 0 5 0
1 189 0 5 0
1 195 0 5 0
1 201 0 5 0
1 207 0 2 0
1 210 0 8 0
1 219 0 8 0
1 228 0 8 0
1 237 0 8 0
1 246 0 8 0
1 255 0 3 0
1 259 0 1 0
1 260 0 1 0
1 261 0 5 0
1 267 0 1 0
1 268 0 1 0
0 269 6 1 4 2 9 14 18
0 270 6 2 4 3 27 15 19
0 273 7 2 3 30 37 43
0 276 7 2 3 4 28 52
0 279 6 1 4 5 10 53 20
0 280 6 3 4 6 11 16 56
0 284 6 1 4 60 44 69 72
0 285 6 1 2 31 70
0 286 6 1 3 61 71 74
0 287 7 2 3 32 76 81
0 290 7 1 3 33 77 45
0 291 7 1 3 34 38 82
0 292 7 1 3 35 39 46
0 293 7 1 3 62 78 83
0 294 7 1 3 63 79 47
0 295 7 1 3 64 40 84
0 296 7 1 3 65 41 48
0 297 7 1 2 85 86
0 298 3 2 2 87 88
0 301 6 1 2 92 97
0 302 3 1 2 93 98
0 303 6 1 2 102 107
0 304 3 1 2 103 108
0 305 6 1 2 112 117
0 306 3 1 2 113 118
0 307 6 1 2 122 127
0 308 3 1 2 123 128
0 309 7 1 2 12 139
0 310 5 5 1 268
0 316 7 1 2 54 140
0 317 7 1 2 21 141
0 318 7 1 2 152 142
0 319 6 2 2 66 157
0 322 4 1 2 22 49
0 323 7 1 2 23 50
0 324 6 1 2 160 166
0 325 3 1 2 161 167
0 326 6 1 2 172 178
0 327 3 1 2 173 179
0 328 6 1 2 184 190
0 329 3 1 2 185 191
0 330 6 1 2 196 202
0 331 3 1 2 197 203
0 332 7 1 2 211 94
0 333 7 1 2 212 99
0 334 7 1 2 213 104
0 335 7 1 2 214 109
0 336 7 1 2 215 114
0 337 7 1 2 256 259
0 338 7 1 2 216 119
0 339 7 1 2 257 260
0 340 7 1 2 217 124
0 341 7 1 2 258 267
0 342 5 1 1 269
0 343 5 1 1 274
0 344 3 1 2 271 275
0 345 5 1 1 277
0 346 5 1 1 278
0 347 5 1 1 279
0 348 4 1 2 281 284
0 349 3 1 2 282 285
0 350 3 1 2 283 286
0 351 5 1 1 293
0 352 5 1 1 294
0 353 5 1 1 295
0 354 5 1 1 296
0 355 6 1 2 89 299
0 356 7 1 2 90 300
0 357 6 2 2 301 302
0 360 6 2 2 303 304
0 363 6 2 2 305 306
0 366 6 2 2 307 308
0 369 5 5 1 311
0 375 4 1 2 322 323
0 376 6 2 2 324 325
0 379 6 2 2 326 327
0 382 6 2 2 328 329
0 385 6 2 2 330 331
3 388 9 0 1 290
3 389 9 0 1 291
3 390 9 0 1 292
3 391 9 0 1 297
0 392 3 1 2 272 343
0 393 5 5 1 345
0 399 5 1 1 346
0 400 7 1 2 348 73
0 401 5 1 1 349
0 402 5 1 1 350
0 403 5 1 1 355
0 404 5 1 1 358
0 405 5 1 1 361
0 406 7 1 2 359 362
0 407 5 1 1 364
0 408 5 1 1 367
0 409 7 1 2 365 368
0 410 6 1 2 347 352
0 411 5 1 1 377
0 412 5 1 1 380
0 413 7 1 2 378 381
0 414 5 1 1 383
0 415 5 1 1 386
0 416 7 1 2 384 387
0 417 7 1 2 218 370
3 418 9 0 1 342
3 419 9 0 1 344
3 420 9 0 1 351
3 421 9 0 1 353
3 422 9 0 1 354
3 423 9 0 1 356
0 424 5 1 1 400
0 425 7 1 2 404 405
0 426 7 1 2 407 408
0 427 7 4 3 320 394 57
0 432 7 4 3 395 24 288
0 437 6 4 3 396 289 58
0 442 6 1 4 375 67 158 397
0 443 6 1 3 398 321 25
0 444 7 1 2 411 412
0 445 7 1 2 414 415
3 446 9 0 1 392
3 447 9 0 1 399
3 448 9 0 1 401
3 449 9 0 1 402
3 450 9 0 1 403
0 451 5 8 1 424
0 460 4 2 2 406 425
0 463 4 2 2 409 426
0 466 6 8 2 442 410
0 475 7 1 2 144 428
0 476 7 1 2 312 433
0 477 7 1 2 147 429
0 478 7 1 2 313 434
0 479 7 1 2 150 430
0 480 7 1 2 314 435
0 481 7 1 2 154 431
0 482 7 1 2 315 436
0 483 6 4 2 443 7
0 488 3 1 2 371 438
0 489 3 1 2 372 439
0 490 3 1 2 373 440
0 491 3 1 2 374 441
0 492 4 2 2 413 444
0 495 4 2 2 416 445
0 498 6 1 2 131 461
0 499 3 1 2 132 462
0 500 6 1 2 464 136
0 501 3 1 2 465 137
0 502 7 1 2 95 467
0 503 4 1 2 475 476
0 504 7 1 2 100 468
0 505 4 1 2 477 478
0 506 7 1 2 105 469
0 507 4 1 2 479 480
0 508 7 1 2 110 470
0 509 4 1 2 481 482
0 510 7 1 2 145 484
0 511 7 1 2 115 471
0 512 7 1 2 148 485
0 513 7 1 2 120 472
0 514 7 1 2 151 486
0 515 7 1 2 125 473
0 516 7 1 2 155 487
0 517 7 1 2 129 474
0 518 6 1 2 133 493
0 519 3 1 2 134 494
0 520 6 1 2 496 208
0 521 3 1 2 497 209
0 522 7 1 2 452 162
0 523 7 1 2 453 168
0 524 7 1 2 454 174
0 525 7 1 2 455 180
0 526 7 1 2 456 186
0 527 6 1 2 457 192
0 528 6 1 2 458 198
0 529 6 1 2 459 204
0 530 6 2 2 498 499
0 533 6 2 2 500 501
0 536 4 1 2 309 502
0 537 4 1 2 316 504
0 538 4 1 2 317 506
0 539 4 1 2 318 508
0 540 4 1 2 510 511
0 541 4 1 2 512 513
0 542 4 1 2 514 515
0 543 4 1 2 516 517
0 544 6 2 2 518 519
0 547 6 2 2 520 521
0 550 5 1 1 531
0 551 5 1 1 534
0 552 7 1 2 532 535
0 553 6 3 2 536 503
0 557 6 3 2 537 505
0 561 6 3 2 538 507
0 565 6 3 2 539 509
0 569 6 3 2 488 540
0 573 6 3 2 489 541
0 577 6 3 2 490 542
0 581 6 3 2 491 543
0 585 5 1 1 545
0 586 5 1 1 548
0 587 7 1 2 546 549
0 588 7 1 2 550 551
0 589 7 1 2 585 586
0 590 6 2 2 554 163
0 593 3 2 2 555 164
0 596 7 1 2 247 556
0 597 6 2 2 558 169
0 600 3 4 2 559 170
0 605 7 1 2 248 560
0 606 6 2 2 562 175
0 609 3 5 2 563 176
0 615 7 1 2 249 564
0 616 6 2 2 566 181
0 619 3 4 2 567 182
0 624 7 1 2 250 568
0 625 6 2 2 570 187
0 628 3 2 2 571 188
0 631 7 1 2 251 572
0 632 6 2 2 574 193
0 635 3 4 2 575 194
0 640 7 1 2 252 576
0 641 6 2 2 578 199
0 644 3 5 2 579 200
0 650 7 1 2 253 580
0 651 6 2 2 582 205
0 654 3 4 2 583 206
0 659 7 1 2 254 584
0 660 4 1 2 552 588
0 661 4 1 2 587 589
0 662 5 2 1 591
0 665 7 3 2 594 592
0 669 4 1 2 596 522
0 670 5 2 1 598
0 673 7 3 2 601 599
0 677 4 1 2 605 523
0 678 5 3 1 607
0 682 7 3 2 610 608
0 686 4 1 2 615 524
0 687 5 4 1 617
0 692 7 3 2 620 618
0 696 4 1 2 624 525
0 697 5 2 1 626
0 700 7 3 2 629 627
0 704 4 1 2 631 526
0 705 5 2 1 633
0 708 7 3 2 636 634
0 712 4 1 2 337 640
0 713 5 3 1 642
0 717 7 3 2 645 643
0 721 4 1 2 339 650
0 722 5 4 1 652
0 727 7 3 2 655 653
0 731 4 1 2 341 659
0 732 6 1 2 656 262
0 733 6 1 3 646 657 263
0 734 6 1 4 637 647 658 264
0 735 5 1 1 663
0 736 7 1 2 229 666
0 737 7 1 2 238 664
0 738 5 1 1 671
0 739 7 1 2 230 674
0 740 7 1 2 239 672
0 741 5 1 1 679
0 742 7 1 2 231 683
0 743 7 1 2 240 680
0 744 5 1 1 688
0 745 7 1 2 232 693
0 746 7 1 2 241 689
0 747 5 1 1 698
0 748 7 1 2 233 701
0 749 7 1 2 242 699
0 750 5 1 1 706
0 751 7 1 2 234 709
0 752 7 1 2 243 707
0 753 5 1 1 714
0 754 7 1 2 235 718
0 755 7 1 2 244 715
0 756 5 1 1 723
0 757 4 1 2 728 265
0 758 7 1 2 729 266
0 759 7 1 2 236 730
0 760 7 1 2 245 724
0 761 6 1 2 648 725
0 762 6 1 2 638 716
0 763 6 1 3 639 649 726
0 764 6 1 2 611 690
0 765 6 1 2 602 681
0 766 6 1 3 603 612 691
3 767 9 0 1 660
3 768 9 0 1 661
0 769 4 1 2 736 737
0 770 4 1 2 739 740
0 771 4 1 2 742 743
0 772 4 1 2 745 746
0 773 6 3 4 750 762 763 734
0 777 4 1 2 748 749
0 778 6 2 3 753 761 733
0 781 4 1 2 751 752
0 782 6 2 2 756 732
0 785 4 1 2 754 755
0 786 4 1 2 757 758
0 787 4 1 2 759 760
0 788 4 1 2 702 774
0 789 7 1 2 703 775
0 790 4 1 2 710 779
0 791 7 1 2 711 780
0 792 4 1 2 719 783
0 793 7 1 2 720 784
0 794 7 1 2 220 786
0 795 6 1 2 630 776
0 796 6 5 2 795 747
0 802 4 1 2 788 789
0 803 4 1 2 790 791
0 804 4 1 2 792 793
0 805 4 1 2 340 794
0 806 4 1 2 694 797
0 807 7 1 2 695 798
0 808 7 1 2 221 802
0 809 7 1 2 222 803
0 810 7 1 2 223 804
0 811 6 1 4 805 787 731 529
0 812 6 1 2 621 799
0 813 6 1 3 613 622 800
0 814 6 1 4 604 614 623 801
0 815 6 3 4 738 765 766 814
0 819 6 2 3 741 764 813
0 822 6 2 2 744 812
0 825 4 1 2 806 807
0 826 4 1 2 335 808
0 827 4 1 2 336 809
0 828 4 1 2 338 810
0 829 5 1 1 811
0 830 4 1 2 667 816
0 831 7 1 2 668 817
0 832 4 1 2 675 820
0 833 7 1 2 676 821
0 834 4 1 2 684 823
0 835 7 1 2 685 824
0 836 7 1 2 224 825
0 837 6 1 3 826 777 704
0 838 6 1 4 827 781 712 527
0 839 6 1 4 828 785 721 528
0 840 5 1 1 829
0 841 6 1 2 818 595
0 842 4 1 2 830 831
0 843 4 1 2 832 833
0 844 4 1 2 834 835
0 845 4 1 2 334 836
0 846 5 1 1 837
0 847 5 1 1 838
0 848 5 1 1 839
0 849 7 1 2 735 841
3 850 9 0 1 840
0 851 7 1 2 225 842
0 852 7 1 2 226 843
0 853 7 1 2 227 844
0 854 6 1 3 845 772 696
0 855 5 1 1 846
0 856 5 1 1 847
0 857 5 1 1 848
0 858 5 1 1 849
0 859 4 1 2 417 851
0 860 4 1 2 332 852
0 861 4 1 2 333 853
0 862 5 1 1 854
3 863 9 0 1 855
3 864 9 0 1 856
3 865 9 0 1 857
3 866 9 0 1 858
0 867 6 1 3 859 769 669
0 868 6 1 3 860 770 677
0 869 6 1 3 861 771 686
0 870 5 1 1 862
0 871 5 1 1 867
0 872 5 1 1 868
0 873 5 1 1 869
3 874 9 0 1 870
0 875 5 1 1 871
0 876 5 1 1 872
0 877 5 1 1 873
3 878 9 0 1 875
3 879 9 0 1 876
3 880 9 0 1 877
2 2 1 1
2 3 1 1
2 4 1 1
2 5 1 1
2 6 1 1
2 7 1 1
2 9 1 8
2 10 1 8
2 11 1 8
2 12 1 8
2 14 1 13
2 15 1 13
2 16 1 13
2 18 1 17
2 19 1 17
2 20 1 17
2 21 1 17
2 22 1 17
2 23 1 17
2 24 1 17
2 25 1 17
2 27 1 26
2 28 1 26
2 30 1 29
2 31 1 29
2 32 1 29
2 33 1 29
2 34 1 29
2 35 1 29
2 37 1 36
2 38 1 36
2 39 1 36
2 40 1 36
2 41 1 36
2 43 1 42
2 44 1 42
2 45 1 42
2 46 1 42
2 47 1 42
2 48 1 42
2 49 1 42
2 50 1 42
2 52 1 51
2 53 1 51
2 54 1 51
2 56 1 55
2 57 1 55
2 58 1 55
2 60 1 59
2 61 1 59
2 62 1 59
2 63 1 59
2 64 1 59
2 65 1 59
2 66 1 59
2 67 1 59
2 69 1 68
2 70 1 68
2 71 1 68
2 76 1 75
2 77 1 75
2 78 1 75
2 79 1 75
2 81 1 80
2 82 1 80
2 83 1 80
2 84 1 80
2 92 1 91
2 93 1 91
2 94 1 91
2 95 1 91
2 97 1 96
2 98 1 96
2 99 1 96
2 100 1 96
2 102 1 101
2 103 1 101
2 104 1 101
2 105 1 101
2 107 1 106
2 108 1 106
2 109 1 106
2 110 1 106
2 112 1 111
2 113 1 111
2 114 1 111
2 115 1 111
2 117 1 116
2 118 1 116
2 119 1 116
2 120 1 116
2 122 1 121
2 123 1 121
2 124 1 121
2 125 1 121
2 127 1 126
2 128 1 126
2 129 1 126
2 131 1 130
2 132 1 130
2 133 1 130
2 134 1 130
2 136 1 135
2 137 1 135
2 139 1 138
2 140 1 138
2 141 1 138
2 142 1 138
2 144 1 143
2 145 1 143
2 147 1 146
2 148 1 146
2 150 1 149
2 151 1 149
2 154 1 153
2 155 1 153
2 157 1 156
2 158 1 156
2 160 1 159
2 161 1 159
2 162 1 159
2 163 1 159
2 164 1 159
2 166 1 165
2 167 1 165
2 168 1 165
2 169 1 165
2 170 1 165
2 172 1 171
2 173 1 171
2 174 1 171
2 175 1 171
2 176 1 171
2 178 1 177
2 179 1 177
2 180 1 177
2 181 1 177
2 182 1 177
2 184 1 183
2 185 1 183
2 186 1 183
2 187 1 183
2 188 1 183
2 190 1 189
2 191 1 189
2 192 1 189
2 193 1 189
2 194 1 189
2 196 1 195
2 197 1 195
2 198 1 195
2 199 1 195
2 200 1 195
2 202 1 201
2 203 1 201
2 204 1 201
2 205 1 201
2 206 1 201
2 208 1 207
2 209 1 207
2 211 1 210
2 212 1 210
2 213 1 210
2 214 1 210
2 215 1 210
2 216 1 210
2 217 1 210
2 218 1 210
2 220 1 219
2 221 1 219
2 222 1 219
2 223 1 219
2 224 1 219
2 225 1 219
2 226 1 219
2 227 1 219
2 229 1 228
2 230 1 228
2 231 1 228
2 232 1 228
2 233 1 228
2 234 1 228
2 235 1 228
2 236 1 228
2 238 1 237
2 239 1 237
2 240 1 237
2 241 1 237
2 242 1 237
2 243 1 237
2 244 1 237
2 245 1 237
2 247 1 246
2 248 1 246
2 249 1 246
2 250 1 246
2 251 1 246
2 252 1 246
2 253 1 246
2 254 1 246
2 256 1 255
2 257 1 255
2 258 1 255
2 262 1 261
2 263 1 261
2 264 1 261
2 265 1 261
2 266 1 261
2 271 1 270
2 272 1 270
2 274 1 273
2 275 1 273
2 277 1 276
2 278 1 276
2 281 1 280
2 282 1 280
2 283 1 280
2 288 1 287
2 289 1 287
2 299 1 298
2 300 1 298
2 311 1 310
2 312 1 310
2 313 1 310
2 314 1 310
2 315 1 310
2 320 1 319
2 321 1 319
2 358 1 357
2 359 1 357
2 361 1 360
2 362 1 360
2 364 1 363
2 365 1 363
2 367 1 366
2 368 1 366
2 370 1 369
2 371 1 369
2 372 1 369
2 373 1 369
2 374 1 369
2 377 1 376
2 378 1 376
2 380 1 379
2 381 1 379
2 383 1 382
2 384 1 382
2 386 1 385
2 387 1 385
2 394 1 393
2 395 1 393
2 396 1 393
2 397 1 393
2 398 1 393
2 428 1 427
2 429 1 427
2 430 1 427
2 431 1 427
2 433 1 432
2 434 1 432
2 435 1 432
2 436 1 432
2 438 1 437
2 439 1 437
2 440 1 437
2 441 1 437
2 452 1 451
2 453 1 451
2 454 1 451
2 455 1 451
2 456 1 451
2 457 1 451
2 458 1 451
2 459 1 451
2 461 1 460
2 462 1 460
2 464 1 463
2 465 1 463
2 467 1 466
2 468 1 466
2 469 1 466
2 470 1 466
2 471 1 466
2 472 1 466
2 473 1 466
2 474 1 466
2 484 1 483
2 485 1 483
2 486 1 483
2 487 1 483
2 493 1 492
2 494 1 492
2 496 1 495
2 497 1 495
2 531 1 530
2 532 1 530
2 534 1 533
2 535 1 533
2 545 1 544
2 546 1 544
2 548 1 547
2 549 1 547
2 554 1 553
2 555 1 553
2 556 1 553
2 558 1 557
2 559 1 557
2 560 1 557
2 562 1 561
2 563 1 561
2 564 1 561
2 566 1 565
2 567 1 565
2 568 1 565
2 570 1 569
2 571 1 569
2 572 1 569
2 574 1 573
2 575 1 573
2 576 1 573
2 578 1 577
2 579 1 577
2 580 1 577
2 582 1 581
2 583 1 581
2 584 1 581
2 591 1 590
2 592 1 590
2 594 1 593
2 595 1 593
2 598 1 597
2 599 1 597
2 601 1 600
2 602 1 600
2 603 1 600
2 604 1 600
2 607 1 606
2 608 1 606
2 610 1 609
2 611 1 609
2 612 1 609
2 613 1 609
2 614 1 609
2 617 1 616
2 618 1 616
2 620 1 619
2 621 1 619
2 622 1 619
2 623 1 619
2 626 1 625
2 627 1 625
2 629 1 628
2 630 1 628
2 633 1 632
2 634 1 632
2 636 1 635
2 637 1 635
2 638 1 635
2 639 1 635
2 642 1 641
2 643 1 641
2 645 1 644
2 646 1 644
2 647 1 644
2 648 1 644
2 649 1 644
2 652 1 651
2 653 1 651
2 655 1 654
2 656 1 654
2 657 1 654
2 658 1 654
2 663 1 662
2 664 1 662
2 666 1 665
2 667 1 665
2 668 1 665
2 671 1 670
2 672 1 670
2 674 1 673
2 675 1 673
2 676 1 673
2 679 1 678
2 680 1 678
2 681 1 678
2 683 1 682
2 684 1 682
2 685 1 682
2 688 1 687
2 689 1 687
2 690 1 687
2 691 1 687
2 693 1 692
2 694 1 692
2 695 1 692
2 698 1 697
2 699 1 697
2 701 1 700
2 702 1 700
2 703 1 700
2 706 1 705
2 707 1 705
2 709 1 708
2 710 1 708
2 711 1 708
2 714 1 713
2 715 1 713
2 716 1 713
2 718 1 717
2 719 1 717
2 720 1 717
2 723 1 722
2 724 1 722
2 725 1 722
2 726 1 722
2 728 1 727
2 729 1 727
2 730 1 727
2 774 1 773
2 775 1 773
2 776 1 773
2 779 1 778
2 780 1 778
2 783 1 782
2 784 1 782
2 797 1 796
2 798 1 796
2 799 1 796
2 800 1 796
2 801 1 796
2 816 1 815
2 817 1 815
2 818 1 815
2 820 1 819
2 821 1 819
2 823 1 822
2 824 1 822
