1 1 0 2 0
1 2 0 2 0
1 3 0 2 0
2 4 1 1
2 5 1 2
2 6 1 1
2 7 1 2
0 8 6 2 2 4 5
2 9 1 8
2 10 1 8
2 11 1 10
0 12 6 1 2 6 9
0 13 6 1 2 11 7
0 14 6 2 2 12 13
2 15 1 14
2 16 1 14
2 17 1 3
2 18 1 3
0 19 6 2 2 16 17
2 20 1 19
2 21 1 19
2 22 1 21
2 23 1 21
2 24 1 10
0 25 6 1 2 15 20
0 26 6 1 2 22 18
3 27 6 0 2 25 26
3 28 6 0 2 23 24
