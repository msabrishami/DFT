1 1 0 3 0
1 5 0 3 0
1 9 0 2 0
1 12 0 2 0
1 15 0 2 0
1 18 0 4 0
1 23 0 2 0
1 26 0 2 0
1 29 0 2 0
1 32 0 2 0
1 35 0 2 0
1 38 0 2 0
1 41 0 2 0
1 44 0 2 0
1 47 0 2 0
1 50 0 2 0
1 53 0 1 0
1 54 0 1 0
1 55 0 1 0
1 56 0 1 0
1 57 0 1 0
1 58 0 1 0
1 59 0 1 0
1 60 0 1 0
1 61 0 1 0
1 62 0 1 0
1 63 0 1 0
1 64 0 1 0
1 65 0 1 0
1 66 0 2 0
1 69 0 1 0
1 70 0 2 0
1 73 0 1 0
1 74 0 1 0
1 75 0 1 0
1 76 0 1 0
1 77 0 1 0
1 78 0 1 0
1 79 0 1 0
1 80 0 1 0
1 81 0 1 0
1 82 0 1 0
1 83 0 1 0
1 84 0 1 0
1 85 0 1 0
1 86 0 1 0
1 87 0 1 0
1 88 0 1 0
1 89 0 4 0
1 94 0 2 0
1 97 0 2 0
1 100 0 2 0
1 103 0 2 0
1 106 0 2 0
1 109 0 1 0
1 110 0 1 0
1 111 0 1 0
1 112 0 1 0
1 113 0 1 0
1 114 0 1 0
1 115 0 2 0
1 118 0 2 0
1 121 0 2 0
1 124 0 2 0
1 127 0 2 0
1 130 0 2 0
1 133 0 1 0
1 134 0 1 0
1 135 0 2 0
1 138 0 2 0
1 141 0 2 0
1 144 0 2 0
1 147 0 2 0
1 150 0 1 0
1 151 0 1 0
1 152 0 1 0
1 153 0 1 0
1 154 0 1 0
1 155 0 1 0
1 156 0 1 0
1 157 0 1 0
1 158 0 1 0
1 159 0 1 0
1 160 0 1 0
1 161 0 1 0
1 162 0 1 0
1 163 0 1 0
1 164 0 1 0
1 165 0 1 0
1 166 0 1 0
1 167 0 1 0
1 168 0 1 0
1 169 0 1 0
1 170 0 1 0
1 171 0 1 0
1 172 0 1 0
1 173 0 1 0
1 174 0 1 0
1 175 0 1 0
1 176 0 1 0
1 177 0 1 0
1 178 0 1 0
1 179 0 1 0
1 180 0 1 0
1 181 0 1 0
1 182 0 1 0
1 183 0 1 0
1 184 0 1 0
1 185 0 1 0
1 186 0 1 0
1 187 0 1 0
1 188 0 1 0
1 189 0 1 0
1 190 0 1 0
1 191 0 1 0
1 192 0 1 0
1 193 0 1 0
1 194 0 1 0
1 195 0 1 0
1 196 0 1 0
1 197 0 1 0
1 198 0 1 0
1 199 0 1 0
1 200 0 1 0
1 201 0 1 0
1 202 0 1 0
1 203 0 1 0
1 204 0 1 0
1 205 0 1 0
1 206 0 1 0
1 207 0 1 0
1 208 0 1 0
1 209 0 1 0
1 210 0 1 0
1 211 0 1 0
1 212 0 1 0
1 213 0 1 0
1 214 0 1 0
1 215 0 1 0
1 216 0 1 0
1 217 0 1 0
1 218 0 1 0
1 219 0 1 0
1 220 0 1 0
1 221 0 1 0
1 222 0 1 0
1 223 0 1 0
1 224 0 1 0
1 225 0 1 0
1 226 0 1 0
1 227 0 1 0
1 228 0 1 0
1 229 0 1 0
1 230 0 1 0
1 231 0 1 0
1 232 0 1 0
1 233 0 1 0
1 234 0 1 0
1 235 0 1 0
1 236 0 1 0
1 237 0 1 0
1 238 0 1 0
1 239 0 1 0
1 240 0 1 0
3 241 0 0 0 
1 242 0 2 0
1 245 0 2 0
1 248 0 2 0
1 251 0 2 0
1 254 0 2 0
1 257 0 2 0
1 260 0 2 0
1 263 0 3 0
1 267 0 3 0
1 271 0 2 0
1 274 0 2 0
1 277 0 2 0
1 280 0 2 0
1 283 0 2 0
1 286 0 2 0
1 289 0 3 0
1 293 0 2 0
1 296 0 2 0
1 299 0 3 0
1 303 0 3 0
1 307 0 2 0
1 310 0 2 0
1 313 0 2 0
1 316 0 2 0
1 319 0 2 0
1 322 0 2 0
1 325 0 2 0
1 328 0 2 0
1 331 0 2 0
1 334 0 2 0
1 337 0 2 0
1 340 0 2 0
1 343 0 2 0
1 346 0 2 0
1 349 0 2 0
1 352 0 2 0
1 355 0 2 0
1 358 0 2 0
1 361 0 2 0
1 364 0 2 0
1 367 0 14 0
1 382 0 4 0
3 387 1 0 1 2
3 388 1 0 1 3
0 467 5 1 1 57
0 469 7 2 2 134 133
3 478 1 0 1 249
3 482 1 0 1 255
3 484 1 0 1 258
3 486 1 0 1 261
3 489 1 0 1 264
3 492 1 0 1 268
0 494 7 2 4 162 172 188 199
3 501 1 0 1 275
3 505 1 0 1 281
3 507 1 0 1 284
3 509 1 0 1 287
3 511 1 0 1 290
3 513 1 0 1 294
3 515 1 0 1 297
3 517 1 0 1 300
3 519 1 0 1 304
0 528 7 2 4 150 184 228 240
3 535 1 0 1 308
3 537 1 0 1 311
3 539 1 0 1 314
3 541 1 0 1 317
3 543 1 0 1 320
3 545 1 0 1 323
3 547 1 0 1 326
3 549 1 0 1 329
3 551 1 0 1 332
3 553 1 0 1 335
3 556 1 0 1 338
3 559 1 0 1 344
3 561 1 0 1 347
3 563 1 0 1 350
3 565 1 0 1 353
3 567 1 0 1 356
3 569 1 0 1 359
3 571 1 0 1 362
3 573 1 0 1 365
0 575 7 2 4 183 182 185 186
0 578 7 2 4 210 152 218 230
3 582 5 0 1 16
0 585 5 1 1 6
0 590 1 2 1 4
0 593 5 2 1 7
0 596 5 2 1 8
0 599 5 4 1 291
0 604 5 4 1 301
0 609 5 4 1 305
0 614 1 10 1 39
0 625 1 2 1 17
0 628 6 3 2 13 10
0 632 6 3 2 14 11
0 636 1 4 1 40
0 641 5 1 1 246
0 642 5 1 1 250
3 643 1 0 1 252
0 644 5 6 1 253
0 651 5 5 1 256
0 657 1 2 1 107
0 660 5 5 1 259
0 666 5 5 1 262
0 672 5 1 1 265
0 673 5 1 1 269
0 674 5 1 1 108
0 676 1 5 1 19
0 682 1 5 1 20
0 688 7 1 2 383 266
0 689 1 5 1 21
0 695 5 4 1 22
0 700 6 4 2 384 270
0 705 5 1 1 272
0 706 5 1 1 276
3 707 1 0 1 278
0 708 5 6 1 279
0 715 5 5 1 282
0 721 5 5 1 285
0 727 5 5 1 288
0 733 5 1 1 292
0 734 5 7 1 295
0 742 5 5 1 298
0 748 5 1 1 302
0 749 5 1 1 306
0 750 1 4 1 368
0 758 5 1 1 309
0 759 5 2 1 312
0 762 5 5 1 315
0 768 5 5 1 318
0 774 5 5 1 321
0 780 5 5 1 324
0 786 5 7 1 327
0 794 5 5 1 330
0 800 5 5 1 333
0 806 5 5 1 336
0 812 5 1 1 339
3 813 1 0 1 341
0 814 5 6 1 342
0 821 5 5 1 345
0 827 5 5 1 348
0 833 5 5 1 351
0 839 5 5 1 354
0 845 5 7 1 357
0 853 5 5 1 360
0 859 5 5 1 363
0 865 5 5 1 366
0 871 1 2 1 369
3 881 6 0 2 467 585
3 882 5 0 1 393
3 883 5 0 1 397
3 884 5 0 1 395
3 885 5 0 1 391
0 886 7 1 2 394 398
0 887 7 1 2 396 392
3 889 1 0 1 399
3 945 1 0 1 450
0 957 5 6 1 688
0 1028 7 1 2 385 641
0 1029 6 2 2 386 705
0 1109 7 1 2 389 403
3 1110 6 0 2 243 401
3 1111 5 0 1 427
3 1112 6 0 2 244 402
3 1113 6 0 2 390 404
3 1114 5 0 1 428
0 1115 5 1 1 679
0 1116 1 2 1 400
0 1119 1 5 1 429
0 1125 1 6 1 468
0 1132 1 3 1 430
0 1136 1 4 1 470
0 1141 1 5 1 431
0 1147 1 6 1 471
0 1154 1 5 1 432
0 1160 1 6 1 462
0 1167 7 4 2 487 417
0 1174 7 1 2 488 418
0 1175 1 6 1 472
0 1182 1 6 1 463
0 1189 5 4 1 451
0 1194 5 4 1 464
0 1199 5 2 1 473
0 1206 5 4 1 474
0 1211 1 6 1 480
0 1218 5 3 1 540
0 1222 5 2 1 1028
0 1227 1 5 1 433
0 1233 1 6 1 465
0 1240 1 3 1 434
0 1244 1 4 1 466
0 1249 1 6 1 475
0 1256 1 6 1 476
0 1263 1 6 1 481
0 1270 1 6 1 477
0 1277 1 6 1 479
0 1284 1 2 1 490
0 1287 1 2 1 419
0 1290 1 2 1 457
0 1293 1 2 1 452
0 1296 1 2 1 445
0 1299 1 2 1 420
0 1302 1 2 1 439
0 1305 1 2 1 491
0 1308 1 2 1 421
0 1311 1 2 1 422
0 1314 1 2 1 458
0 1317 1 2 1 453
0 1320 1 2 1 446
0 1323 1 2 1 440
0 1326 1 2 1 413
0 1329 1 2 1 409
0 1332 1 2 1 532
0 1335 1 2 1 405
0 1338 1 2 1 518
0 1341 1 2 1 508
0 1344 1 2 1 500
0 1347 1 2 1 524
0 1350 1 2 1 493
0 1353 1 2 1 414
0 1356 1 2 1 410
0 1359 1 2 1 533
0 1362 1 2 1 525
0 1365 1 2 1 406
0 1368 1 2 1 520
0 1371 1 2 1 510
0 1374 1 2 1 502
0 1377 1 2 1 495
0 1380 1 2 1 608
0 1383 1 2 1 602
0 1386 1 2 1 595
0 1389 1 2 1 586
0 1392 1 2 1 579
0 1395 1 2 1 570
0 1398 1 2 1 560
0 1401 1 2 1 552
0 1404 1 2 1 610
0 1407 1 2 1 603
0 1410 1 2 1 597
0 1413 1 2 1 580
0 1416 1 2 1 572
0 1419 1 2 1 562
0 1422 1 2 1 554
0 1425 1 2 1 587
0 1428 1 2 1 435
0 1431 1 2 1 436
0 1434 1 2 1 670
0 1437 1 2 1 664
0 1440 1 2 1 658
0 1443 1 2 1 649
0 1446 1 2 1 640
0 1449 1 2 1 634
0 1452 1 2 1 627
0 1455 1 2 1 621
0 1458 1 2 1 615
0 1461 1 2 1 671
0 1464 1 2 1 665
0 1467 1 2 1 659
0 1470 1 2 1 645
0 1473 1 2 1 635
0 1476 1 2 1 629
0 1479 1 2 1 622
0 1482 1 2 1 650
0 1485 1 2 1 616
3 1489 5 0 1 1109
3 1490 1 0 1 692
0 1537 7 5 2 681 423
0 1551 7 2 2 424 683
0 1649 7 1 2 690 437
0 1703 1 2 1 684
0 1708 4 2 2 685 425
0 1713 1 2 1 686
0 1721 4 2 2 426 687
0 1758 1 2 1 691
3 1781 7 0 2 163 693
0 1782 7 1 2 170 701
0 1783 5 5 1 702
0 1789 5 3 1 714
0 1793 7 1 2 169 703
0 1794 7 1 2 168 704
0 1795 7 1 2 167 709
0 1796 7 1 2 166 716
0 1797 7 1 2 165 717
0 1798 7 1 2 164 718
0 1799 5 5 1 725
0 1805 5 5 1 739
0 1811 7 1 2 177 726
0 1812 7 1 2 176 728
0 1813 7 1 2 175 729
0 1814 7 1 2 174 730
0 1815 7 1 2 173 731
0 1816 7 1 2 157 740
0 1817 7 1 2 156 741
0 1818 7 1 2 155 743
0 1819 7 1 2 154 744
0 1820 7 1 2 153 745
0 1821 5 1 1 857
0 1822 5 1 1 860
0 1828 5 1 1 862
0 1829 5 1 1 864
0 1830 5 1 1 867
0 1832 5 1 1 869
0 1833 5 1 1 872
0 1834 5 1 1 874
0 1835 5 1 1 876
0 1839 5 1 1 878
0 1840 5 1 1 880
0 1841 5 1 1 890
0 1842 5 1 1 892
0 1843 5 1 1 894
0 1845 5 5 1 753
0 1851 5 5 1 761
0 1857 7 1 2 181 754
0 1858 7 1 2 171 755
0 1859 7 1 2 180 756
0 1860 7 1 2 179 757
0 1861 7 1 2 178 760
0 1862 7 1 2 161 763
0 1863 7 1 2 151 764
0 1864 7 1 2 160 765
0 1865 7 1 2 159 766
0 1866 7 1 2 158 767
0 1867 5 1 1 896
0 1868 5 1 1 898
0 1869 5 1 1 900
0 1870 5 1 1 902
0 1871 5 1 1 904
0 1872 5 1 1 906
0 1873 5 1 1 908
0 1874 5 1 1 910
0 1875 5 1 1 912
0 1876 5 1 1 914
0 1877 5 1 1 916
0 1878 5 1 1 918
0 1879 5 1 1 920
0 1880 5 1 1 922
0 1881 5 1 1 924
0 1882 5 1 1 926
0 1883 5 1 1 928
0 1884 5 1 1 930
0 1885 1 6 1 778
0 1892 1 6 1 773
0 1899 1 6 1 779
0 1906 1 6 1 775
0 1913 5 5 1 785
0 1919 1 6 1 776
0 1926 7 1 2 45 787
0 1927 7 1 2 42 788
0 1928 7 1 2 30 789
0 1929 7 1 2 27 790
0 1930 7 1 2 24 791
0 1931 5 1 1 932
0 1932 5 1 1 934
0 1933 5 1 1 936
0 1934 5 1 1 938
0 1935 5 1 1 940
0 1936 5 1 1 942
0 1937 5 1 1 944
0 1938 5 1 1 947
0 1939 5 1 1 949
0 1940 5 1 1 951
0 1941 5 1 1 953
0 1942 5 1 1 955
0 1943 5 1 1 958
0 1944 5 1 1 960
0 1945 5 1 1 962
0 1946 5 1 1 964
0 1947 5 5 1 804
0 1953 5 3 1 817
0 1957 7 1 2 209 805
0 1958 7 1 2 216 807
0 1959 7 1 2 215 808
0 1960 7 1 2 214 809
0 1961 7 1 2 213 818
0 1962 7 1 2 212 819
0 1963 7 1 2 211 820
0 1965 5 1 1 966
0 1966 7 1 2 796 438
0 1967 5 1 1 968
0 1968 5 1 1 970
0 1969 5 1 1 972
0 1970 5 1 1 974
0 1971 5 1 1 976
0 1972 5 1 1 978
0 1973 5 1 1 980
0 1974 5 1 1 982
0 1975 5 1 1 984
0 1976 5 1 1 986
0 1977 5 5 1 822
0 1983 5 5 1 829
0 1989 7 1 2 642 823
0 1990 7 1 2 441 824
0 1991 7 1 2 447 825
0 1992 7 1 2 674 826
0 1993 7 1 2 454 828
0 1994 7 1 2 459 830
0 1995 7 1 2 672 831
0 1996 7 1 2 673 832
0 1997 5 5 1 836
0 2003 1 6 1 777
0 2010 7 1 2 48 837
0 2011 7 1 2 36 838
0 2012 7 1 2 33 840
0 2013 7 1 2 51 841
0 2014 7 1 2 67 842
0 2015 5 1 1 988
0 2016 5 1 1 990
0 2017 5 1 1 992
0 2018 5 1 1 994
0 2019 5 1 1 996
0 2020 5 1 1 998
0 2021 5 1 1 1000
0 2022 5 1 1 1002
0 2023 5 1 1 1004
0 2024 1 6 1 781
0 2031 1 6 1 782
0 2038 1 6 1 783
0 2045 1 6 1 784
0 2052 5 5 1 843
0 2058 5 5 1 850
0 2064 7 1 2 706 844
0 2065 7 1 2 496 846
0 2066 7 1 2 503 847
0 2067 7 1 2 512 848
0 2068 7 1 2 521 849
0 2069 7 1 2 733 851
0 2070 7 1 2 526 852
0 2071 7 1 2 534 854
0 2072 7 1 2 748 855
0 2073 7 1 2 749 856
0 2074 1 2 1 769
0 2081 1 2 1 770
0 2086 1 2 1 797
0 2107 6 1 2 861 1821
0 2108 6 1 2 858 1822
0 2110 5 1 1 1013
0 2111 6 1 2 1014 1832
0 2112 6 1 2 877 1834
0 2113 6 1 2 875 1835
0 2114 5 1 1 1017
0 2115 6 1 2 1018 1839
0 2117 5 1 1 1019
0 2171 5 1 1 1021
0 2172 6 1 2 1022 1965
0 2230 5 1 1 1015
0 2231 1 2 1 1006
0 2235 1 2 1 1011
0 2239 3 1 2 1023 1782
0 2240 3 1 2 1024 710
0 2241 3 1 2 1025 1793
0 2242 3 1 2 1026 1794
0 2243 3 1 2 1027 1795
0 2244 3 1 2 1030 1796
0 2245 3 1 2 1031 1797
0 2246 3 1 2 1032 1798
0 2247 3 1 2 1033 1811
0 2248 3 1 2 1034 1812
0 2249 3 1 2 1035 1813
0 2250 3 1 2 1036 1814
0 2251 3 1 2 1037 1815
0 2252 3 1 2 1038 1816
0 2253 3 1 2 1039 1817
0 2254 3 1 2 1040 1818
0 2255 3 1 2 1041 1819
0 2256 3 1 2 1042 1820
0 2257 6 9 2 2107 2108
0 2267 5 1 1 1168
0 2268 6 1 2 870 2110
0 2269 6 4 2 2112 2113
0 2274 6 1 2 879 2114
0 2275 5 1 1 1170
0 2277 7 1 2 142 1043
0 2278 7 1 2 148 1044
0 2279 7 1 2 139 1045
0 2280 7 1 2 145 1046
0 2281 7 1 2 136 1047
0 2282 7 1 2 143 1048
0 2283 7 1 2 149 1049
0 2284 7 1 2 140 1050
0 2285 7 1 2 146 1051
0 2286 7 1 2 137 1052
0 2287 5 5 1 1053
0 2293 5 5 1 1059
0 2299 7 1 2 104 1054
0 2300 7 1 2 131 1055
0 2301 7 1 2 128 1056
0 2302 7 1 2 125 1057
0 2303 7 1 2 101 1058
0 2304 7 1 2 105 1060
0 2305 7 1 2 132 1061
0 2306 7 1 2 129 1062
0 2307 7 1 2 126 1063
0 2308 7 1 2 102 1064
0 2309 5 5 1 1065
0 2315 5 5 1 1071
0 2321 7 1 2 116 1066
0 2322 7 1 2 119 1067
0 2323 7 1 2 98 1068
0 2324 7 1 2 95 1069
0 2325 7 1 2 122 1070
0 2326 7 1 2 117 1072
0 2327 7 1 2 120 1073
0 2328 7 1 2 99 1074
0 2329 7 1 2 96 1075
0 2330 7 1 2 123 1076
0 2331 5 5 1 1082
0 2337 7 1 2 208 1077
0 2338 7 1 2 198 1078
0 2339 7 1 2 207 1079
0 2340 7 1 2 206 1080
0 2341 7 1 2 205 1081
0 2342 7 1 2 46 1083
0 2343 7 1 2 43 1084
0 2344 7 1 2 31 1085
0 2345 7 1 2 28 1086
0 2346 7 1 2 25 1087
0 2347 3 1 2 1088 810
0 2348 3 1 2 1089 1957
0 2349 3 1 2 1090 1958
0 2350 3 1 2 1091 1959
0 2351 3 1 2 1092 1960
0 2352 3 1 2 1093 1961
0 2353 3 1 2 1094 1962
0 2354 3 1 2 1095 1963
0 2355 6 1 2 967 2171
0 2356 5 1 1 1172
0 2357 6 1 2 1173 1967
0 2358 7 1 2 114 1096
0 2359 7 1 2 113 1097
0 2360 7 1 2 111 1098
0 2361 7 1 2 87 1099
0 2362 7 1 2 112 1100
0 2363 7 1 2 88 1101
0 2364 7 1 2 247 1102
0 2365 7 1 2 273 1103
0 2366 7 1 2 548 1104
0 2367 7 1 2 71 1105
0 2368 5 5 1 1120
0 2374 7 1 2 193 1106
0 2375 7 1 2 192 1107
0 2376 7 1 2 191 1108
0 2377 7 1 2 190 1117
0 2378 7 1 2 189 1118
0 2379 7 1 2 49 1121
0 2380 7 1 2 37 1122
0 2381 7 1 2 34 1123
0 2382 7 1 2 52 1124
0 2383 7 1 2 68 1126
0 2384 5 5 1 1127
0 2390 5 5 1 1134
0 2396 7 1 2 58 1128
0 2397 7 1 2 77 1129
0 2398 7 1 2 78 1130
0 2399 7 1 2 59 1131
0 2400 7 1 2 81 1133
0 2401 7 1 2 80 1135
0 2402 7 1 2 79 1137
0 2403 7 1 2 60 1138
0 2404 7 1 2 61 1139
0 2405 7 1 2 62 1140
0 2406 5 5 1 1142
0 2412 5 5 1 1149
0 2418 7 1 2 69 1143
0 2419 7 1 2 72 1144
0 2420 7 1 2 74 1145
0 2421 7 1 2 76 1146
0 2422 7 1 2 75 1148
0 2423 7 1 2 73 1150
0 2424 7 1 2 53 1151
0 2425 7 1 2 54 1152
0 2426 7 1 2 55 1153
0 2427 7 1 2 56 1155
0 2428 7 1 2 82 1156
0 2429 7 1 2 65 1157
0 2430 7 1 2 83 1158
0 2431 7 1 2 84 1159
0 2432 7 1 2 85 1161
0 2433 7 1 2 64 1162
0 2434 7 1 2 63 1163
0 2435 7 1 2 86 1164
0 2436 7 1 2 109 1165
0 2437 7 1 2 110 1166
0 2441 7 1 2 2239 694
0 2442 7 3 2 2240 696
0 2446 7 3 2 2241 697
0 2450 7 3 2 2242 698
0 2454 7 3 2 2243 699
0 2458 7 3 2 2244 711
0 2462 7 3 2 2247 719
0 2466 7 3 2 2248 720
0 2470 7 3 2 2249 722
0 2474 7 3 2 2250 723
0 2478 7 3 2 2251 724
0 2482 7 5 2 2252 732
0 2488 7 7 2 2253 735
0 2496 7 5 2 2254 736
0 2502 7 5 2 2255 737
0 2508 7 5 2 2256 738
0 2523 6 5 2 2268 2111
0 2533 6 3 2 2274 2115
0 2537 5 1 1 1178
0 2538 3 3 2 2278 1858
0 2542 3 3 2 2279 1859
0 2546 3 3 2 2280 1860
0 2550 3 3 2 2281 1861
0 2554 3 6 2 2283 1863
0 2561 3 5 2 2284 1864
0 2567 3 5 2 2285 1865
0 2573 3 5 2 2286 1866
0 2604 3 2 2 2338 1927
0 2607 3 3 2 2339 1928
0 2611 3 3 2 2340 1929
0 2615 3 3 2 2341 1930
0 2619 7 6 2 2348 798
0 2626 7 5 2 2349 799
0 2632 7 5 2 2350 801
0 2638 7 5 2 2351 802
0 2644 7 5 2 2352 811
0 2650 6 2 2 2355 2172
0 2653 6 1 2 969 2356
0 2654 3 3 2 2359 1990
0 2658 3 3 2 2360 1991
0 2662 3 3 2 2361 1992
0 2666 3 3 2 2362 1993
0 2670 3 3 2 2363 1994
0 2674 3 5 2 2366 834
0 2680 3 2 2 2367 835
0 2688 3 3 2 2374 2010
0 2692 3 3 2 2375 2011
0 2696 3 3 2 2376 2012
0 2700 3 3 2 2377 2013
0 2704 3 3 2 2378 2014
0 2728 7 1 2 2347 803
0 2729 3 3 2 2429 2065
0 2733 3 3 2 2430 2066
0 2737 3 3 2 2431 2067
0 2741 3 3 2 2432 2068
0 2745 3 3 2 2433 2069
0 2749 3 3 2 2434 2070
0 2753 3 3 2 2435 2071
0 2757 3 3 2 2436 2072
0 2761 3 3 2 2437 2073
0 2765 5 1 1 1176
0 2766 7 2 2 2354 815
0 2769 7 2 2 2353 816
0 2772 7 2 2 2246 712
0 2775 7 2 2 2245 713
0 2778 3 2 2 2282 1862
0 2781 3 2 2 2358 1989
0 2784 3 2 2 2365 1996
0 2787 3 2 2 2364 1995
0 2790 3 2 2 2337 1926
0 2793 3 2 2 2277 1857
0 2796 3 2 2 2428 2064
0 2866 7 1 2 1180 1007
0 2867 7 1 2 1181 1008
0 2868 7 1 2 1183 1009
0 2869 7 1 2 1184 1010
0 2878 7 1 2 1191 1012
0 2913 7 1 2 204 1196
0 2914 7 1 2 203 1197
0 2915 7 1 2 202 1198
0 2916 7 1 2 201 1200
0 2917 7 1 2 200 1201
0 2918 7 1 2 235 1202
0 2919 7 1 2 234 1203
0 2920 7 1 2 233 1204
0 2921 7 1 2 232 1205
0 2922 7 1 2 231 1207
0 2923 7 1 2 197 1208
0 2924 7 1 2 187 1209
0 2925 7 1 2 196 1210
0 2926 7 1 2 195 1212
0 2927 7 1 2 194 1213
0 2928 7 1 2 227 1214
0 2929 7 1 2 217 1215
0 2930 7 1 2 226 1216
0 2931 7 1 2 225 1217
0 2932 7 1 2 224 1219
0 2933 7 1 2 239 1220
0 2934 7 1 2 229 1221
0 2935 7 1 2 238 1223
0 2936 7 1 2 237 1224
0 2937 7 1 2 236 1225
0 2988 6 1 2 2653 2357
0 3005 7 1 2 223 1226
0 3006 7 1 2 222 1228
0 3007 7 1 2 221 1229
0 3008 7 1 2 220 1230
0 3009 7 1 2 219 1231
0 3020 7 1 2 812 1232
0 3021 7 1 2 617 1234
0 3022 7 1 2 623 1235
0 3023 7 1 2 630 1236
0 3024 7 1 2 637 1237
0 3025 7 1 2 646 1238
0 3026 7 1 2 652 1239
0 3027 7 1 2 661 1241
0 3028 7 1 2 667 1242
0 3029 7 1 2 675 1243
0 3032 7 1 2 758 1245
0 3033 7 1 2 550 1246
0 3034 7 1 2 555 1247
0 3035 7 1 2 564 1248
0 3036 7 1 2 574 1250
0 3037 7 1 2 581 1251
0 3038 7 1 2 588 1252
0 3039 7 1 2 598 1253
0 3040 7 1 2 605 1254
0 3041 7 1 2 611 1255
0 3061 1 2 1 1185
0 3064 1 2 1 1186
0 3067 1 2 1 1192
0 3070 1 2 1 1193
0 3073 5 2 1 2728
0 3080 5 2 1 2441
0 3096 7 1 2 460 1444
0 3097 7 3 2 455 1436
0 3101 7 5 2 771 1429
0 3107 7 6 2 448 1421
0 3114 7 7 2 442 1412
0 3122 7 3 2 1334 1187
0 3126 3 3 2 746 2866
0 3130 7 1 2 1336 1188
0 3131 3 2 2 747 2869
0 3134 7 1 2 1337 1190
0 3135 5 1 1 1342
0 3136 7 1 2 461 1445
0 3137 7 2 2 456 1438
0 3140 7 3 2 772 1430
0 3144 7 4 2 449 1423
0 3149 7 5 2 443 1414
0 3155 7 3 2 1343 1195
0 3159 3 3 2 1174 2878
0 3167 5 1 1 1540
0 3168 7 1 2 415 1327
0 3169 7 3 2 411 1319
0 3173 7 4 2 536 1312
0 3178 7 5 2 527 1301
0 3184 7 1 2 407 1294
0 3185 7 3 2 522 1388
0 3189 7 5 2 514 1381
0 3195 7 6 2 504 1373
0 3202 7 7 2 497 1364
0 3210 7 1 2 416 1328
0 3211 7 3 2 412 1321
0 3215 7 5 2 538 1313
0 3221 7 6 2 1303 529
0 3228 7 1 2 408 1295
0 3229 7 2 2 523 1390
0 3232 7 3 2 516 1382
0 3236 7 4 2 506 1375
0 3241 7 5 2 498 1366
0 3247 3 3 2 2913 2299
0 3251 3 3 2 2914 2300
0 3255 3 3 2 2915 2301
0 3259 3 3 2 2916 2302
0 3263 3 3 2 2917 2303
0 3267 3 5 2 2918 2304
0 3273 3 7 2 2919 2305
0 3281 3 5 2 2920 2306
0 3287 3 5 2 2921 2307
0 3293 3 5 2 2922 2308
0 3299 3 3 2 2924 2322
0 3303 3 3 2 2925 2323
0 3307 3 3 2 2926 2324
0 3311 3 3 2 2927 2325
0 3315 3 6 2 2929 2327
0 3322 3 5 2 2930 2328
0 3328 3 5 2 2931 2329
0 3334 3 5 2 2932 2330
0 3340 3 2 2 2934 2343
0 3343 3 5 2 2935 2344
0 3349 3 5 2 2936 2345
0 3355 3 5 2 2937 2346
0 3361 7 1 2 1528 1289
0 3362 7 1 2 1525 1285
0 3363 7 1 2 1522 1281
0 3364 7 1 2 1519 1278
0 3365 7 1 2 1516 1274
0 3366 7 1 2 1513 1360
0 3367 7 1 2 1510 1355
0 3368 7 1 2 1507 1351
0 3369 7 1 2 1504 1346
0 3370 7 1 2 1472 1271
0 3371 7 1 2 1468 1267
0 3372 7 1 2 1463 1264
0 3373 7 1 2 1459 1260
0 3374 7 1 2 1454 1257
0 3375 7 3 2 2988 1451
0 3379 7 1 2 1453 1966
0 3380 5 1 1 1542
0 3381 7 2 2 483 1396
0 3384 3 5 2 3005 2379
0 3390 3 7 2 3006 2380
0 3398 3 5 2 3007 2381
0 3404 3 5 2 3008 2382
0 3410 3 5 2 3009 2383
0 3416 3 3 2 3021 2397
0 3420 3 3 2 3022 2398
0 3424 3 3 2 3023 2399
0 3428 3 3 2 3024 2400
0 3432 3 3 2 3025 2401
0 3436 3 3 2 3026 2402
0 3440 3 3 2 3027 2403
0 3444 3 3 2 3028 2404
0 3448 3 3 2 3029 2405
0 3452 5 1 1 1548
0 3453 5 1 1 1550
0 3454 3 3 2 3034 2420
0 3458 3 3 2 3035 2421
0 3462 3 3 2 3036 2422
0 3466 3 3 2 3037 2423
0 3470 3 3 2 3038 2424
0 3474 3 3 2 3039 2425
0 3478 3 3 2 3040 2426
0 3482 3 3 2 3041 2427
0 3486 5 1 1 1553
0 3487 1 2 1 1447
0 3490 1 2 1 1439
0 3493 1 2 1 1432
0 3496 1 2 1 1424
0 3499 1 2 1 1415
0 3502 1 2 1 1339
0 3507 4 2 2 751 2868
0 3510 1 2 1 1340
0 3515 4 2 2 444 1417
0 3518 1 2 1 1448
0 3521 1 2 1 1441
0 3524 1 2 1 1433
0 3527 1 2 1 1426
0 3530 1 2 1 1418
0 3535 1 2 1 1420
0 3539 1 2 1 1435
0 3542 1 2 1 1427
0 3545 1 2 1 1450
0 3548 1 2 1 1442
0 3551 5 1 1 1531
0 3552 5 1 1 1533
0 3553 1 2 1 1258
0 3557 1 2 1 1265
0 3560 1 2 1 1261
0 3563 1 2 1 1272
0 3566 1 2 1 1268
0 3569 5 1 1 1535
0 3570 5 1 1 1538
0 3571 1 2 1 1367
0 3574 1 2 1 1384
0 3577 1 2 1 1376
0 3580 1 2 1 1297
0 3583 1 2 1 1391
0 3586 1 2 1 1315
0 3589 1 2 1 1304
0 3592 1 2 1 1330
0 3595 1 2 1 1322
0 3598 1 2 1 1331
0 3601 1 2 1 1324
0 3604 1 2 1 1316
0 3607 1 2 1 1298
0 3610 1 2 1 1393
0 3613 1 2 1 1385
0 3616 1 2 1 1378
0 3619 1 2 1 1306
0 3622 1 2 1 1369
0 3625 4 2 2 530 1307
0 3628 4 2 2 499 1370
0 3631 1 2 1 1333
0 3634 1 2 1 1325
0 3637 1 2 1 1318
0 3640 1 2 1 1309
0 3643 1 2 1 1300
0 3646 1 2 1 1394
0 3649 1 2 1 1387
0 3652 1 2 1 1379
0 3655 1 2 1 1372
0 3658 4 2 2 1310 531
0 3661 1 2 1 1477
0 3664 1 2 1 1478
0 3667 1 2 1 1529
0 3670 1 2 1 1291
0 3673 1 2 1 1526
0 3676 1 2 1 1286
0 3679 1 2 1 1523
0 3682 1 2 1 1282
0 3685 1 2 1 1517
0 3688 1 2 1 1275
0 3691 1 2 1 1514
0 3694 1 2 1 1361
0 3697 1 2 1 1511
0 3700 1 2 1 1357
0 3703 1 2 1 1508
0 3706 1 2 1 1352
0 3709 1 2 1 1520
0 3712 1 2 1 1279
0 3715 1 2 1 1505
0 3718 1 2 1 1348
0 3721 1 2 1 1501
0 3724 1 2 1 1498
0 3727 1 2 1 1495
0 3730 1 2 1 1487
0 3733 1 2 1 1492
0 3736 1 2 1 1474
0 3739 1 2 1 1273
0 3742 1 2 1 1469
0 3745 1 2 1 1269
0 3748 1 2 1 1465
0 3751 1 2 1 1266
0 3754 1 2 1 1460
0 3757 1 2 1 1262
0 3760 1 2 1 1456
0 3763 1 2 1 1259
0 3766 1 2 1 1457
0 3769 1 2 1 1466
0 3772 1 2 1 1462
0 3775 1 2 1 1475
0 3778 1 2 1 1471
0 3781 5 1 1 1544
0 3782 5 1 1 1546
0 3783 3 2 2 2928 2326
0 3786 3 2 2 2933 2342
0 3789 3 2 2 2923 2321
0 3792 1 2 1 1488
0 3795 1 2 1 1496
0 3798 1 2 1 1493
0 3801 1 2 1 1502
0 3804 1 2 1 1499
0 3807 1 2 1 1397
0 3810 1 2 1 1403
0 3813 1 2 1 1399
0 3816 1 2 1 1408
0 3819 1 2 1 1349
0 3822 1 2 1 1358
0 3825 1 2 1 1354
0 3828 1 2 1 1276
0 3831 1 2 1 1363
0 3834 1 2 1 1283
0 3837 1 2 1 1280
0 3840 1 2 1 1292
0 3843 1 2 1 1288
0 3846 1 2 1 1409
0 3849 1 2 1 1405
0 3852 1 2 1 1400
0 3855 1 2 1 1484
0 3858 1 2 1 1506
0 3861 1 2 1 1512
0 3864 1 2 1 1509
0 3867 1 2 1 1518
0 3870 1 2 1 1515
0 3873 1 2 1 1524
0 3876 1 2 1 1521
0 3879 1 2 1 1530
0 3882 1 2 1 1527
0 3885 3 2 2 3033 2419
0 3888 3 2 2 3032 2418
0 3891 3 2 2 3020 2396
0 3953 6 1 2 1559 2117
0 3954 5 1 1 1560
0 3955 6 1 2 1561 2537
0 3956 5 1 1 1562
0 3958 5 1 1 1563
0 3964 5 1 1 1565
0 4193 3 3 2 1649 3379
0 4303 3 2 3 752 2867 3130
0 4308 5 1 1 1555
0 4313 5 1 1 1557
0 4326 6 1 2 1534 3551
0 4327 6 1 2 1532 3552
0 4333 6 1 2 1539 3569
0 4334 6 1 2 1536 3570
0 4411 6 1 2 1547 3781
0 4412 6 1 2 1545 3782
0 4463 6 1 2 1952 1828
0 4464 5 1 1 1954
0 4465 6 1 2 1955 1829
0 4466 5 1 1 1956
0 4467 6 1 2 1964 2267
0 4468 5 1 1 1978
0 4469 6 1 2 1979 1830
0 4470 5 1 1 1980
0 4471 6 1 2 1981 1833
0 4472 5 1 1 1982
0 4473 5 1 1 1588
0 4474 5 1 1 1591
0 4475 6 1 2 2001 1840
0 4476 5 1 1 2002
0 4477 6 1 2 2004 1841
0 4478 5 1 1 2005
0 4479 6 1 2 2006 2275
0 4480 5 1 1 2007
0 4481 6 1 2 2008 1842
0 4482 5 1 1 2009
0 4483 6 1 2 2025 1843
0 4484 5 1 1 2026
0 4485 5 1 1 1610
0 4486 5 1 1 1613
0 4487 6 1 2 1020 3954
0 4488 6 1 2 1179 3956
0 4489 5 1 1 2027
0 4490 6 1 2 2028 3958
0 4491 5 1 1 2029
0 4492 5 1 1 2032
0 4493 5 1 1 2034
0 4494 5 1 1 2036
0 4495 5 1 1 2039
0 4496 6 1 2 2040 3964
0 4497 5 1 1 2041
0 4498 5 1 1 2043
0 4499 5 1 1 2046
0 4500 5 1 1 2048
0 4501 5 1 1 2050
0 4502 6 1 2 2051 3167
0 4503 5 1 1 2053
0 4504 5 1 1 2055
0 4505 5 1 1 2057
0 4506 5 1 1 2060
0 4507 6 1 2 2082 1867
0 4508 5 1 1 2083
0 4509 6 1 2 2084 1868
0 4510 5 1 1 2085
0 4511 6 1 2 2087 1869
0 4512 5 1 1 2088
0 4513 6 1 2 2089 1870
0 4514 5 1 1 2090
0 4515 6 1 2 2091 1871
0 4516 5 1 1 2092
0 4517 6 1 2 2093 1872
0 4518 5 1 1 2094
0 4519 6 1 2 2095 1873
0 4520 5 1 1 2096
0 4521 6 1 2 2097 1874
0 4522 5 1 1 2098
0 4523 6 1 2 2099 1875
0 4524 5 1 1 2100
0 4525 6 1 2 2105 1876
0 4526 5 1 1 2106
0 4527 6 1 2 2109 1877
0 4528 5 1 1 2116
0 4529 6 1 2 2118 1878
0 4530 5 1 1 2119
0 4531 6 1 2 2120 1879
0 4532 5 1 1 2121
0 4533 6 1 2 2122 1880
0 4534 5 1 1 2123
0 4535 6 1 2 2124 1881
0 4536 5 1 1 2125
0 4537 6 1 2 2126 1882
0 4538 5 1 1 2127
0 4539 6 1 2 2128 1883
0 4540 5 1 1 2129
0 4541 6 1 2 2130 1884
0 4542 5 1 1 2131
0 4543 5 1 1 2132
0 4544 7 1 2 612 1718
0 4545 7 3 2 606 1712
0 4549 7 5 2 600 1706
0 4555 7 6 2 1698 589
0 4562 7 1 2 583 1693
0 4563 7 2 2 576 1770
0 4566 7 3 2 566 1765
0 4570 7 4 2 557 1760
0 4575 5 1 1 2134
0 4576 7 1 2 613 1719
0 4577 7 3 2 607 1714
0 4581 7 4 2 601 1707
0 4586 7 5 2 591 1699
0 4592 7 1 2 584 1694
0 4593 7 3 2 577 1771
0 4597 7 5 2 568 1766
0 4603 7 6 2 558 1761
0 4610 5 1 1 2136
0 4611 5 1 1 2138
0 4612 5 1 1 2140
0 4613 5 1 1 2142
0 4614 5 1 1 2144
0 4615 5 1 1 2146
0 4616 5 1 1 2148
0 4617 5 1 1 2150
0 4618 5 1 1 2152
0 4619 5 1 1 2154
0 4620 5 1 1 2156
0 4621 5 1 1 2158
0 4622 5 1 1 2160
0 4623 5 1 1 2162
0 4624 5 1 1 2164
0 4625 5 1 1 2166
0 4626 5 1 1 2168
0 4627 5 1 1 2170
0 4628 5 1 1 2174
0 4629 5 1 1 2176
0 4630 7 1 2 1900 1503
0 4631 5 1 1 2178
0 4632 7 1 2 1896 1500
0 4633 5 1 1 2180
0 4634 7 1 2 1893 1497
0 4635 7 1 2 1889 1494
0 4636 5 1 1 2182
0 4637 7 1 2 1886 1491
0 4638 7 1 2 1854 1733
0 4639 7 1 2 1850 1730
0 4640 7 1 2 1847 1727
0 4641 7 1 2 1838 1724
0 4642 5 1 1 2184
0 4643 5 1 1 2186
0 4644 5 1 1 2188
0 4645 5 1 1 2190
0 4646 5 1 1 2192
0 4647 5 1 1 2194
0 4648 5 1 1 2196
0 4649 5 1 1 2198
0 4650 5 1 1 2200
0 4651 5 1 1 2202
0 4652 5 1 1 2204
0 4653 5 1 1 1775
0 4656 7 1 2 677 1826
0 4657 7 3 2 668 1809
0 4661 7 5 2 662 1803
0 4667 7 6 2 1788 653
0 4674 7 1 2 647 1780
0 4675 7 2 2 638 1752
0 4678 7 3 2 631 1747
0 4682 7 4 2 624 1742
0 4687 7 5 2 618 1736
0 4693 5 1 1 2206
0 4694 6 1 2 2207 3380
0 4695 5 1 1 2208
0 4696 5 1 1 2210
0 4697 5 1 1 2212
0 4698 5 1 1 2214
0 4699 5 1 1 2216
0 4700 5 1 1 2218
0 4701 7 1 2 678 1827
0 4702 7 3 2 669 1810
0 4706 7 4 2 663 1804
0 4711 7 5 2 654 1790
0 4717 7 1 2 648 1784
0 4718 7 3 2 639 1753
0 4722 7 5 2 633 1748
0 4728 7 6 2 626 1743
0 4735 7 7 2 619 1737
0 4743 5 1 1 2220
0 4744 5 1 1 2222
0 4745 5 1 1 2234
0 4746 6 1 2 2236 3452
0 4747 5 1 1 2237
0 4748 5 1 1 2258
0 4749 5 1 1 2260
0 4750 5 1 1 2262
0 4751 6 1 2 2263 3453
0 4752 5 1 1 2264
0 4753 5 1 1 2266
0 4754 5 1 1 2271
0 4755 5 1 1 2273
0 4756 7 1 2 1949 1690
0 4757 7 1 2 1924 1687
0 4758 7 1 2 1921 1684
0 4759 7 1 2 1917 1681
0 4760 7 1 2 1914 1678
0 4761 5 1 1 2297
0 4762 7 1 2 1910 1411
0 4763 5 1 1 2310
0 4764 7 1 2 1907 1406
0 4765 5 1 1 2312
0 4766 7 1 2 1903 1402
0 4767 7 1 2 1486 1778
0 4768 5 1 1 2314
0 4769 7 5 2 1757 485
0 4775 5 1 1 2317
0 4776 6 1 2 2318 3486
0 4777 5 1 1 2319
0 4778 5 1 1 2332
0 4779 5 1 1 2334
0 4780 5 1 1 2336
0 4781 5 1 1 2389
0 4782 5 1 1 2392
0 4783 5 1 1 2394
0 4784 3 2 2 1594 3134
0 4789 5 1 1 1984
0 4790 5 2 1 1595
0 4793 5 1 1 1986
0 4794 5 1 1 1988
0 4795 5 1 1 1999
0 4796 1 2 1 1581
0 4799 5 1 1 2062
0 4800 5 1 1 2075
0 4801 5 1 1 2077
0 4802 5 1 1 2079
0 4803 6 2 2 4326 4327
0 4806 6 2 2 4333 4334
0 4809 5 1 1 2101
0 4810 1 2 1 1623
0 4813 5 1 1 2103
0 4814 1 2 1 1642
0 4817 1 2 1 1658
0 4820 1 2 1 1720
0 4823 1 2 1 1715
0 4826 1 2 1 1709
0 4829 1 2 1 1700
0 4832 1 2 1 1695
0 4835 1 2 1 1772
0 4838 1 2 1 1767
0 4841 1 2 1 1762
0 4844 4 2 2 1701 592
0 4847 1 2 1 1722
0 4850 1 2 1 1716
0 4853 1 2 1 1710
0 4856 1 2 1 1696
0 4859 1 2 1 1773
0 4862 1 2 1 1768
0 4865 1 2 1 1763
0 4868 1 2 1 1702
0 4871 4 2 2 594 1704
0 4874 1 2 1 1901
0 4877 1 2 1 1897
0 4880 1 2 1 1894
0 4883 1 2 1 1887
0 4886 1 2 1 1855
0 4889 1 2 1 1734
0 4892 1 2 1 1852
0 4895 1 2 1 1731
0 4898 1 2 1 1848
0 4901 1 2 1 1728
0 4904 1 2 1 1890
0 4907 1 2 1 1844
0 4910 1 2 1 1725
0 4913 1 2 1 1831
0 4916 1 2 1 1823
0 4919 1 2 1 1806
0 4922 1 2 1 1791
0 4925 1 2 1 1785
0 4928 1 2 1 1754
0 4931 1 2 1 1749
0 4934 1 2 1 1744
0 4937 1 2 1 1738
0 4940 4 2 2 1792 655
0 4943 1 2 1 1739
0 4946 1 2 1 1750
0 4949 1 2 1 1745
0 4952 1 2 1 1786
0 4955 1 2 1 1755
0 4958 1 2 1 1807
0 4961 1 2 1 1800
0 4964 1 2 1 1836
0 4967 1 2 1 1824
0 4970 1 2 1 1759
0 4973 1 2 1 1769
0 4976 1 2 1 1764
0 4979 1 2 1 1697
0 4982 1 2 1 1774
0 4985 1 2 1 1711
0 4988 1 2 1 1705
0 4991 1 2 1 1723
0 4994 1 2 1 1717
0 4997 6 2 2 4411 4412
0 5000 1 2 1 1837
0 5003 1 2 1 1825
0 5006 1 2 1 1808
0 5009 1 2 1 1787
0 5012 1 2 1 1756
0 5015 1 2 1 1751
0 5018 1 2 1 1746
0 5021 1 2 1 1801
0 5024 1 2 1 1740
0 5027 4 2 2 656 1802
0 5030 4 2 2 620 1741
0 5033 1 2 1 1726
0 5036 1 2 1 1732
0 5039 1 2 1 1729
0 5042 1 2 1 1735
0 5045 5 1 1 2224
0 5046 5 1 1 2226
0 5047 5 1 1 2228
0 5048 5 1 1 2232
0 5049 1 2 1 1679
0 5052 1 2 1 1685
0 5055 1 2 1 1682
0 5058 1 2 1 1691
0 5061 1 2 1 1688
0 5064 5 1 1 2288
0 5065 5 1 1 2290
0 5066 5 1 1 2292
0 5067 5 1 1 2295
0 5068 1 2 1 1950
0 5071 1 2 1 1692
0 5074 1 2 1 1925
0 5077 1 2 1 1689
0 5080 1 2 1 1922
0 5083 1 2 1 1686
0 5086 1 2 1 1915
0 5089 1 2 1 1680
0 5092 1 2 1 1911
0 5095 1 2 1 1908
0 5098 1 2 1 1904
0 5101 1 2 1 1918
0 5104 1 2 1 1683
0 5107 1 2 1 1779
0 5110 5 1 1 2370
0 5111 5 1 1 2372
0 5112 5 1 1 2385
0 5113 5 1 1 2387
0 5114 1 2 1 1909
0 5117 1 2 1 1905
0 5120 1 2 1 1916
0 5123 1 2 1 1912
0 5126 1 2 1 1923
0 5129 1 2 1 1920
0 5132 1 2 1 1951
0 5135 1 2 1 1948
0 5138 1 2 1 1846
0 5141 1 2 1 1853
0 5144 1 2 1 1849
0 5147 1 2 1 1888
0 5150 1 2 1 1856
0 5153 1 2 1 1895
0 5156 1 2 1 1891
0 5159 1 2 1 1902
0 5162 1 2 1 1898
0 5165 6 1 2 4486 4485
0 5166 6 1 2 4474 4473
0 5167 6 1 2 863 4464
0 5168 6 1 2 866 4466
0 5169 6 1 2 1169 4468
0 5170 6 1 2 868 4470
0 5171 6 1 2 873 4472
0 5172 6 1 2 888 4476
0 5173 6 1 2 891 4478
0 5174 6 1 2 1171 4480
0 5175 6 1 2 893 4482
0 5176 6 1 2 895 4484
0 5177 6 1 2 3953 4487
0 5178 6 1 2 3955 4488
0 5179 6 1 2 1564 4489
0 5180 6 1 2 2033 4491
0 5181 6 1 2 2030 4492
0 5182 6 1 2 2037 4493
0 5183 6 1 2 2035 4494
0 5184 6 1 2 1566 4495
0 5185 6 1 2 2044 4497
0 5186 6 1 2 2042 4498
0 5187 6 1 2 2049 4499
0 5188 6 1 2 2047 4500
0 5189 6 1 2 1541 4501
0 5190 6 1 2 2056 4503
0 5191 6 1 2 2054 4504
0 5192 6 1 2 2061 4505
0 5193 6 1 2 2059 4506
0 5196 6 1 2 897 4508
0 5197 6 1 2 899 4510
0 5198 6 1 2 901 4512
0 5199 6 1 2 903 4514
0 5200 6 1 2 905 4516
0 5201 6 1 2 907 4518
0 5202 6 1 2 909 4520
0 5203 6 1 2 911 4522
0 5204 6 1 2 913 4524
0 5205 6 1 2 915 4526
0 5206 6 1 2 917 4528
0 5207 6 1 2 919 4530
0 5208 6 1 2 921 4532
0 5209 6 1 2 923 4534
0 5210 6 1 2 925 4536
0 5211 6 1 2 927 4538
0 5212 6 1 2 929 4540
0 5213 6 1 2 931 4542
0 5283 6 1 2 2141 4611
0 5284 6 1 2 2139 4612
0 5285 6 1 2 2145 4613
0 5286 6 1 2 2143 4614
0 5287 6 1 2 2149 4615
0 5288 6 1 2 2147 4616
0 5289 6 1 2 2153 4617
0 5290 6 1 2 2151 4618
0 5291 6 1 2 2157 4619
0 5292 6 1 2 2155 4620
0 5293 6 1 2 2161 4621
0 5294 6 1 2 2159 4622
0 5295 6 1 2 2165 4623
0 5296 6 1 2 2163 4624
0 5297 6 1 2 2169 4625
0 5298 6 1 2 2167 4626
0 5299 6 1 2 2175 4627
0 5300 6 1 2 2173 4628
0 5314 6 1 2 2189 4643
0 5315 6 1 2 2187 4644
0 5316 6 1 2 2193 4645
0 5317 6 1 2 2191 4646
0 5318 6 1 2 2197 4647
0 5319 6 1 2 2195 4648
0 5320 6 1 2 2201 4649
0 5321 6 1 2 2199 4650
0 5322 6 1 2 2205 4651
0 5323 6 1 2 2203 4652
0 5324 5 1 1 2407
0 5363 6 1 2 1543 4693
0 5364 6 1 2 2211 4695
0 5365 6 1 2 2209 4696
0 5366 6 1 2 2215 4697
0 5367 6 1 2 2213 4698
0 5425 6 1 2 1549 4745
0 5426 6 1 2 2259 4747
0 5427 6 1 2 2238 4748
0 5429 6 1 2 1552 4750
0 5430 6 1 2 2270 4752
0 5431 6 1 2 2265 4753
0 5432 6 1 2 2276 4754
0 5433 6 1 2 2272 4755
0 5451 6 1 2 1554 4775
0 5452 6 1 2 2333 4777
0 5453 6 1 2 2320 4778
0 5454 6 1 2 2369 4779
0 5455 6 1 2 2335 4780
0 5456 6 1 2 2393 4781
0 5457 6 1 2 2391 4782
0 5469 5 1 1 2410
0 5474 6 1 2 2076 4799
0 5475 6 1 2 2063 4800
0 5476 6 1 2 2080 4801
0 5477 6 1 2 2078 4802
0 5571 6 1 2 2227 5045
0 5572 6 1 2 2225 5046
0 5573 6 1 2 2233 5047
0 5574 6 1 2 2229 5048
0 5584 6 1 2 2291 5064
0 5585 6 1 2 2289 5065
0 5586 6 1 2 2296 5066
0 5587 6 1 2 2294 5067
0 5602 6 1 2 2373 5110
0 5603 6 1 2 2371 5111
0 5604 6 1 2 2388 5112
0 5605 6 1 2 2386 5113
0 5631 6 1 2 5324 4653
0 5632 6 7 2 4463 5167
0 5640 6 13 2 4465 5168
0 5654 6 15 2 4467 5169
0 5670 6 12 2 4469 5170
0 5683 6 6 2 4471 5171
0 5690 6 6 2 4475 5172
0 5697 6 9 2 4477 5173
0 5707 6 10 2 4479 5174
0 5718 6 9 2 4481 5175
0 5728 6 6 2 4483 5176
0 5735 5 1 1 5177
0 5736 6 3 2 5179 4490
0 5740 6 3 2 5180 5181
0 5744 6 2 2 5182 5183
0 5747 6 3 2 5184 4496
0 5751 6 3 2 5185 5186
0 5755 6 2 2 5187 5188
0 5758 6 3 2 5189 4502
0 5762 6 3 2 5190 5191
0 5766 6 2 2 5192 5193
0 5769 5 1 1 2581
0 5770 5 1 1 2583
0 5771 6 6 2 4507 5196
0 5778 6 10 2 4509 5197
0 5789 6 9 2 4511 5198
0 5799 6 7 2 4513 5199
0 5807 6 13 2 4515 5200
0 5821 6 15 2 4517 5201
0 5837 6 12 2 4519 5202
0 5850 6 5 2 4521 5203
0 5856 6 6 2 4523 5204
0 5863 6 6 2 4525 5205
0 5870 6 10 2 4527 5206
0 5881 6 10 2 4529 5207
0 5892 6 5 2 4531 5208
0 5898 6 6 2 4533 5209
0 5905 6 9 2 4535 5210
0 5915 6 10 2 4537 5211
0 5926 6 9 2 4539 5212
0 5936 6 6 2 4541 5213
0 5943 5 1 1 2589
0 5944 6 1 2 2591 1931
0 5945 5 1 1 2592
0 5946 6 1 2 2593 1932
0 5947 5 1 1 2594
0 5948 6 1 2 2595 1933
0 5949 5 1 1 2596
0 5950 6 1 2 2597 1934
0 5951 5 1 1 2598
0 5952 6 1 2 2599 1935
0 5953 5 1 1 2600
0 5954 6 1 2 2601 1936
0 5955 5 1 1 2602
0 5956 6 1 2 2603 1937
0 5957 5 1 1 2605
0 5958 6 1 2 2606 1938
0 5959 5 1 1 2608
0 5960 7 5 2 1480 2569
0 5966 5 1 1 2609
0 5967 6 1 2 2612 1939
0 5968 5 1 1 2613
0 5969 6 1 2 2614 1940
0 5970 5 1 1 2616
0 5971 6 1 2 2617 1941
0 5972 5 1 1 2618
0 5973 6 1 2 2620 1942
0 5974 5 1 1 2621
0 5975 6 1 2 2622 1943
0 5976 5 1 1 2623
0 5977 6 1 2 2624 1944
0 5978 5 1 1 2625
0 5979 6 1 2 2627 1945
0 5980 5 1 1 2628
0 5981 7 7 2 1481 2570
0 5989 6 1 2 2629 1946
0 5990 5 1 1 2630
0 5991 6 4 2 5283 5284
0 5996 6 3 2 5285 5286
0 6000 6 2 2 5287 5288
0 6003 6 5 2 5289 5290
0 6009 6 4 2 5291 5292
0 6014 6 3 2 5293 5294
0 6018 6 2 2 5295 5296
0 6021 6 1 2 5297 5298
0 6022 6 1 2 5299 5300
0 6023 5 1 1 2634
0 6024 6 1 2 2635 4629
0 6025 5 1 1 2636
0 6026 6 1 2 2637 4631
0 6027 5 1 1 2639
0 6028 6 1 2 2640 4633
0 6029 5 1 1 2641
0 6030 6 1 2 2642 4636
0 6031 5 1 1 2643
0 6032 5 1 1 2646
0 6033 5 1 1 2648
0 6034 5 1 1 2651
0 6035 5 1 1 2655
0 6036 5 1 1 2657
0 6037 5 1 1 2660
0 6038 6 1 2 2661 4642
0 6039 5 1 1 2663
0 6040 5 1 1 2665
0 6041 6 5 2 5314 5315
0 6047 6 4 2 5316 5317
0 6052 6 3 2 5318 5319
0 6056 6 2 2 5320 5321
0 6059 6 1 2 5322 5323
0 6060 6 1 2 2668 1968
0 6061 5 1 1 2669
0 6062 6 1 2 2671 1969
0 6063 5 1 1 2672
0 6064 6 1 2 2673 1970
0 6065 5 1 1 2675
0 6066 6 1 2 2676 1971
0 6067 5 1 1 2677
0 6068 6 1 2 2678 1972
0 6069 5 1 1 2679
0 6070 6 1 2 2681 1973
0 6071 5 1 1 2682
0 6072 6 1 2 2683 1974
0 6073 5 1 1 2684
0 6074 6 1 2 2685 1975
0 6075 5 1 1 2686
0 6076 6 1 2 2687 1976
0 6077 5 1 1 2689
0 6078 5 1 1 2690
0 6079 6 3 2 5363 4694
0 6083 6 3 2 5364 5365
0 6087 6 2 2 5366 5367
0 6090 5 1 1 2693
0 6091 6 1 2 2694 4699
0 6092 5 1 1 2695
0 6093 5 1 1 2698
0 6094 5 1 1 2701
0 6095 5 1 1 2703
0 6096 5 1 1 2714
0 6097 6 1 2 2715 4700
0 6098 5 1 1 2716
0 6099 5 1 1 2718
0 6100 5 1 1 2720
0 6101 5 1 1 2722
0 6102 5 1 1 2735
0 6103 6 1 2 2738 2015
0 6104 5 1 1 2739
0 6105 6 1 2 2740 2016
0 6106 5 1 1 2742
0 6107 6 1 2 2743 2017
0 6108 5 1 1 2744
0 6109 6 1 2 2746 2018
0 6110 5 1 1 2747
0 6111 6 1 2 2748 2019
0 6112 5 1 1 2750
0 6113 6 1 2 2751 2020
0 6114 5 1 1 2752
0 6115 6 1 2 2754 2021
0 6116 5 1 1 2755
0 6117 6 1 2 2756 2022
0 6118 5 1 1 2758
0 6119 6 1 2 2759 2023
0 6120 5 1 1 2760
0 6121 5 1 1 2768
0 6122 6 1 2 2770 4743
0 6123 5 1 1 2771
0 6124 5 1 1 2774
0 6125 6 1 2 2777 4744
0 6126 5 1 1 2779
0 6127 6 3 2 5425 4746
0 6131 6 3 2 5426 5427
0 6135 5 1 1 2780
0 6136 6 1 2 2782 4749
0 6137 6 3 2 5429 4751
0 6141 6 3 2 5430 5431
0 6145 6 2 2 5432 5433
0 6148 5 1 1 2795
0 6149 5 1 1 2798
0 6150 5 1 1 2800
0 6151 5 1 1 2802
0 6152 5 1 1 2804
0 6153 5 1 1 2806
0 6154 5 1 1 2808
0 6155 5 1 1 2810
0 6156 5 1 1 2812
0 6157 6 1 2 2813 4761
0 6158 5 1 1 2814
0 6159 6 1 2 2815 4763
0 6160 5 1 1 2816
0 6161 6 1 2 2817 4765
0 6162 5 1 1 2818
0 6163 5 1 1 2820
0 6164 6 1 2 2822 4768
0 6165 5 1 1 2823
0 6166 6 3 2 5451 4776
0 6170 6 3 2 5452 5453
0 6174 6 2 2 5454 5455
0 6177 6 3 2 5456 5457
0 6181 5 1 1 2824
0 6182 5 1 1 2826
0 6183 5 1 1 2828
0 6184 5 1 1 2830
0 6185 5 1 1 2840
0 6186 6 1 2 2841 4783
0 6187 5 1 1 2842
0 6188 5 1 1 2844
0 6189 5 1 1 2846
0 6190 5 1 1 2848
0 6191 5 1 1 2575
0 6192 6 1 2 2576 2230
0 6193 5 1 1 2577
0 6194 6 1 2 2578 2765
0 6195 5 1 1 2579
0 6196 6 2 2 5476 5477
0 6199 6 2 2 5474 5475
0 6202 5 1 1 2585
0 6203 5 1 1 2587
0 6204 1 2 1 2571
0 6207 1 2 1 2443
0 6210 1 2 1 2572
0 6213 5 1 1 2631
0 6214 1 2 1 2472
0 6217 4 2 2 1483 2574
0 6220 1 2 1 2505
0 6223 5 1 1 2706
0 6224 5 1 1 2708
0 6225 5 1 1 2710
0 6226 5 1 1 2712
0 6227 5 1 1 2724
0 6228 5 1 1 2726
0 6229 5 1 1 2730
0 6230 5 1 1 2732
0 6231 5 1 1 2762
0 6232 1 2 1 2535
0 6235 5 1 1 2764
0 6236 1 2 1 2560
0 6239 5 1 1 2783
0 6240 5 1 1 2786
0 6241 5 1 1 2789
0 6242 5 1 1 2792
0 6243 6 2 2 5573 5574
0 6246 6 2 2 5571 5572
0 6249 6 2 2 5586 5587
0 6252 6 2 2 5584 5585
0 6255 5 1 1 2832
0 6256 5 1 1 2834
0 6257 5 1 1 2836
0 6258 5 1 1 2838
0 6259 5 1 1 2850
0 6260 5 1 1 2852
0 6261 5 1 1 2854
0 6262 5 1 1 2856
0 6263 6 2 2 5604 5605
0 6266 6 2 2 5602 5603
0 6540 6 1 2 933 5945
0 6541 6 1 2 935 5947
0 6542 6 1 2 937 5949
0 6543 6 1 2 939 5951
0 6544 6 1 2 941 5953
0 6545 6 1 2 943 5955
0 6546 6 1 2 946 5957
0 6547 6 1 2 948 5959
0 6555 6 1 2 950 5968
0 6556 6 1 2 952 5970
0 6557 6 1 2 954 5972
0 6558 6 1 2 956 5974
0 6559 6 1 2 959 5976
0 6560 6 1 2 961 5978
0 6561 6 1 2 963 5980
0 6569 6 1 2 965 5990
0 6594 6 1 2 2177 6023
0 6595 6 1 2 2179 6025
0 6596 6 1 2 2181 6027
0 6597 6 1 2 2183 6029
0 6598 6 1 2 2647 6031
0 6599 6 1 2 2645 6032
0 6600 6 1 2 2652 6033
0 6601 6 1 2 2649 6034
0 6602 6 1 2 2659 6035
0 6603 6 1 2 2656 6036
0 6604 6 1 2 2185 6037
0 6605 6 1 2 2667 6039
0 6606 6 1 2 2664 6040
0 6621 6 1 2 971 6061
0 6622 6 1 2 973 6063
0 6623 6 1 2 975 6065
0 6624 6 1 2 977 6067
0 6625 6 1 2 979 6069
0 6626 6 1 2 981 6071
0 6627 6 1 2 983 6073
0 6628 6 1 2 985 6075
0 6629 6 1 2 987 6077
0 6639 6 1 2 2217 6090
0 6640 6 1 2 2699 6092
0 6641 6 1 2 2697 6093
0 6642 6 1 2 2705 6094
0 6643 6 1 2 2702 6095
0 6644 6 1 2 2219 6096
0 6645 6 1 2 2719 6098
0 6646 6 1 2 2717 6099
0 6647 6 1 2 2723 6100
0 6648 6 1 2 2721 6101
0 6649 6 1 2 989 6104
0 6650 6 1 2 991 6106
0 6651 6 1 2 993 6108
0 6652 6 1 2 995 6110
0 6653 6 1 2 997 6112
0 6654 6 1 2 999 6114
0 6655 6 1 2 1001 6116
0 6656 6 1 2 1003 6118
0 6657 6 1 2 1005 6120
0 6658 6 1 2 2221 6121
0 6659 6 1 2 2776 6123
0 6660 6 1 2 2773 6124
0 6661 6 1 2 2223 6126
0 6668 6 1 2 2261 6135
0 6677 6 1 2 2799 6148
0 6678 6 1 2 2797 6149
0 6679 6 1 2 2803 6150
0 6680 6 1 2 2801 6151
0 6681 6 1 2 2807 6152
0 6682 6 1 2 2805 6153
0 6683 6 1 2 2811 6154
0 6684 6 1 2 2809 6155
0 6685 6 1 2 2298 6156
0 6686 6 1 2 2311 6158
0 6687 6 1 2 2313 6160
0 6688 6 1 2 2821 6162
0 6689 6 1 2 2819 6163
0 6690 6 1 2 2316 6165
0 6702 6 1 2 2827 6181
0 6703 6 1 2 2825 6182
0 6704 6 1 2 2831 6183
0 6705 6 1 2 2829 6184
0 6706 6 1 2 2395 6185
0 6707 6 1 2 2845 6187
0 6708 6 1 2 2843 6188
0 6709 6 1 2 2849 6189
0 6710 6 1 2 2847 6190
0 6711 6 1 2 1016 6191
0 6712 6 1 2 1177 6193
0 6729 6 1 2 2709 6223
0 6730 6 1 2 2707 6224
0 6731 6 1 2 2713 6225
0 6732 6 1 2 2711 6226
0 6733 6 1 2 2727 6227
0 6734 6 1 2 2725 6228
0 6735 6 1 2 2734 6229
0 6736 6 1 2 2731 6230
0 6741 6 1 2 2788 6239
0 6742 6 1 2 2785 6240
0 6743 6 1 2 2794 6241
0 6744 6 1 2 2791 6242
0 6751 6 1 2 2835 6255
0 6752 6 1 2 2833 6256
0 6753 6 1 2 2839 6257
0 6754 6 1 2 2837 6258
0 6755 6 1 2 2853 6259
0 6756 6 1 2 2851 6260
0 6757 6 1 2 2857 6261
0 6758 6 1 2 2855 6262
0 6761 5 1 1 3164
0 6762 7 3 5 2910 2898 2883 2865 2858
0 6766 7 1 2 2859 1567
0 6767 7 1 3 2870 2860 1570
0 6768 7 1 4 2884 2861 1575 2871
0 6769 7 1 5 2899 2885 2862 1582 2872
0 6770 7 1 2 2873 1571
0 6771 7 1 3 2886 1576 2874
0 6772 7 1 4 2900 2887 1583 2875
0 6773 7 1 4 2911 2888 2876 2901
0 6774 7 1 2 2877 1572
0 6775 7 1 3 2889 1577 2879
0 6776 7 1 4 2902 2890 1584 2880
0 6777 7 1 2 2891 1578
0 6778 7 1 3 2903 2892 1585
0 6779 7 1 3 2912 2893 2904
0 6780 7 1 2 2894 1579
0 6781 7 1 3 2905 2895 1586
0 6782 7 1 2 2906 1587
0 6783 7 1 2 2938 2907
0 6784 7 2 5 2947 2975 2956 2941 2966
0 6787 7 1 2 2942 1596
0 6788 7 1 3 2948 2943 1598
0 6789 7 1 4 2957 2944 1601 2949
0 6790 7 1 5 2967 2958 2945 1605 2950
0 6791 7 1 2 2951 1599
0 6792 7 1 3 2959 1602 2952
0 6793 7 1 4 2968 2960 1606 2953
0 6794 7 1 2 1603 2961
0 6795 7 1 3 2969 2962 1607
0 6796 7 1 2 2970 1608
0 6797 5 2 1 2981
0 6800 5 2 1 2984
0 6803 5 2 1 2990
0 6806 5 2 1 2993
0 6809 5 2 1 2998
0 6812 5 2 1 3001
0 6815 1 2 1 2987
0 6818 1 2 1 2989
0 6821 1 2 1 2996
0 6824 1 2 1 2997
0 6827 1 2 1 3004
0 6830 1 2 1 3010
0 6833 7 2 4 3113 3047 3017 3011
0 6836 7 1 2 3012 1616
0 6837 7 1 3 3018 3013 1619
0 6838 7 1 4 3048 3014 1624 3019
0 6839 7 1 2 3030 1620
0 6840 7 1 3 3049 1625 3031
0 6841 7 1 3 3115 3050 3042
0 6842 7 1 2 3043 1621
0 6843 7 1 3 3051 1626 3044
0 6844 7 1 2 3052 1627
0 6845 7 2 5 3119 3099 3082 3065 3056
0 6848 7 1 2 3057 1628
0 6849 7 1 3 3066 3058 1631
0 6850 7 1 4 3083 3059 1636 3068
0 6851 7 1 5 3100 3084 3060 1643 3069
0 6852 7 1 2 3071 1632
0 6853 7 1 3 3085 1637 3072
0 6854 7 1 4 3102 3086 1644 3074
0 6855 7 1 4 3120 3087 3075 3103
0 6856 7 1 2 3076 1633
0 6857 7 1 3 3088 1638 3077
0 6858 7 1 4 3104 3089 1645 3078
0 6859 7 1 2 3090 1639
0 6860 7 1 3 3105 3091 1646
0 6861 7 1 3 3121 3092 3106
0 6862 7 1 2 3093 1640
0 6863 7 1 3 3108 3094 1647
0 6864 7 1 2 3109 1648
0 6865 7 1 2 3116 3053
0 6866 7 1 2 3123 3110
0 6867 7 2 4 3139 3165 3152 3127
0 6870 7 1 2 3128 1650
0 6871 7 1 3 3141 3129 1653
0 6872 7 1 4 3153 3132 1659 3142
0 6873 7 1 2 3143 1654
0 6874 7 1 3 3154 1660 3145
0 6875 7 1 3 3166 3156 3146
0 6876 7 1 2 3147 1655
0 6877 7 1 3 1661 3157 3148
0 6878 7 1 2 3158 1662
0 6879 7 1 2 3170 3160
0 6880 7 1 2 3161 1663
0 6881 7 2 5 3180 3216 3192 3172 3204
0 6884 7 1 2 3174 1664
0 6885 7 1 3 3181 3175 1666
0 6886 7 1 4 3193 3176 1669 3182
0 6887 7 1 5 3205 3194 3177 1673 3183
0 6888 7 1 2 3186 1667
0 6889 7 1 3 3196 1670 3187
0 6890 7 1 4 3206 3197 1674 3188
0 6891 7 1 2 1671 3198
0 6892 7 1 3 3207 3199 1675
0 6893 7 1 2 3208 1676
0 6894 6 6 2 5944 6540
0 6901 6 10 2 5946 6541
0 6912 6 10 2 5948 6542
0 6923 6 5 2 5950 6543
0 6929 6 6 2 5952 6544
0 6936 6 9 2 5954 6545
0 6946 6 10 2 5956 6546
0 6957 6 9 2 5958 6547
0 6967 6 1 2 3331 4575
0 6968 5 1 1 3332
0 6969 5 1 1 3333
0 6970 6 6 2 5967 6555
0 6977 6 10 2 5969 6556
0 6988 6 9 2 5971 6557
0 6998 6 7 2 5973 6558
0 7006 6 13 2 5975 6559
0 7020 6 15 2 5977 6560
0 7036 6 12 2 5979 6561
0 7049 6 5 2 5989 6569
0 7055 6 1 2 3336 4610
0 7056 5 1 1 3337
0 7057 7 2 4 6021 3248 3244 3239
0 7060 7 1 2 3240 3362
0 7061 7 1 3 3245 3242 3363
0 7062 7 1 4 3249 3243 3364 3246
0 7063 7 1 5 6022 3266 3262 3257 3250
0 7064 7 1 2 3252 3366
0 7065 7 1 3 3258 3253 3367
0 7066 7 1 4 3264 3254 3368 3260
0 7067 7 1 5 3268 3265 3256 3369 3261
0 7068 6 4 2 6594 6024
0 7073 6 3 2 6595 6026
0 7077 6 2 2 6596 6028
0 7080 6 5 2 6597 6030
0 7086 6 4 2 6598 6599
0 7091 6 3 2 6600 6601
0 7095 6 2 2 6602 6603
0 7098 6 1 2 6604 6038
0 7099 6 1 2 6605 6606
0 7100 7 2 5 6059 3283 3279 3275 3269
0 7103 7 1 2 3270 3371
0 7104 7 1 3 3276 3271 3372
0 7105 7 1 4 3280 3272 3373 3277
0 7106 7 1 5 3284 3282 3274 3374 3278
0 7107 6 6 2 6060 6621
0 7114 6 10 2 6062 6622
0 7125 6 10 2 6064 6623
0 7136 6 5 2 6066 6624
0 7142 6 6 2 6068 6625
0 7149 6 9 2 6070 6626
0 7159 6 10 2 6072 6627
0 7170 6 9 2 6074 6628
0 7180 6 6 2 6076 6629
0 7187 5 1 1 3344
0 7188 5 2 1 3285
0 7191 5 2 1 3289
0 7194 6 3 2 6639 6091
0 7198 6 3 2 6640 6641
0 7202 6 2 2 6642 6643
0 7205 6 3 2 6644 6097
0 7209 6 3 2 6645 6646
0 7213 6 2 2 6647 6648
0 7216 1 2 1 3292
0 7219 1 2 1 3294
0 7222 6 6 2 6103 6649
0 7229 6 10 2 6105 6650
0 7240 6 9 2 6107 6651
0 7250 6 7 2 6109 6652
0 7258 6 13 2 6111 6653
0 7272 6 15 2 6113 6654
0 7288 6 12 2 6115 6655
0 7301 6 5 2 6117 6656
0 7307 6 6 2 6119 6657
0 7314 6 3 2 6658 6122
0 7318 6 3 2 6659 6660
0 7322 6 2 2 6125 6661
0 7325 5 2 1 3295
0 7328 5 2 1 3298
0 7331 6 2 2 6668 6136
0 7334 5 2 1 3302
0 7337 5 2 1 3306
0 7340 1 2 1 3310
0 7343 1 2 1 3312
0 7346 6 4 2 6677 6678
0 7351 6 3 2 6679 6680
0 7355 6 2 2 6681 6682
0 7358 6 5 2 6683 6684
0 7364 6 4 2 6685 6157
0 7369 6 3 2 6686 6159
0 7373 6 2 2 6687 6161
0 7376 6 1 2 6688 6689
0 7377 6 1 2 6164 6690
0 7378 5 2 1 3313
0 7381 5 2 1 3317
0 7384 5 2 1 3323
0 7387 6 3 2 6702 6703
0 7391 6 2 2 6704 6705
0 7394 6 3 2 6706 6186
0 7398 6 3 2 6707 6708
0 7402 6 2 2 6709 6710
0 7405 1 2 1 3320
0 7408 1 2 1 3321
0 7411 1 2 1 3217
0 7414 1 2 1 3179
0 7417 1 2 1 3190
0 7420 1 2 1 3200
0 7423 1 2 1 3209
0 7426 1 2 1 2976
0 7429 1 2 1 2946
0 7432 1 2 1 2954
0 7435 1 2 1 2963
0 7438 1 2 1 2971
0 7441 6 2 2 6192 6711
0 7444 6 2 2 6194 6712
0 7447 1 2 1 2939
0 7450 1 2 1 2908
0 7453 1 2 1 2863
0 7456 1 2 1 2896
0 7459 1 2 1 2881
0 7462 1 2 1 2882
0 7465 1 2 1 2940
0 7468 1 2 1 2909
0 7471 1 2 1 2864
0 7474 1 2 1 2897
0 7477 5 1 1 3326
0 7478 5 1 1 3329
0 7479 1 2 1 3117
0 7482 1 2 1 3054
0 7485 1 2 1 3015
0 7488 1 2 1 3045
0 7491 1 2 1 3118
0 7494 1 2 1 3055
0 7497 1 2 1 3016
0 7500 1 2 1 3046
0 7503 1 2 1 3124
0 7506 1 2 1 3111
0 7509 1 2 1 3062
0 7512 1 2 1 3095
0 7515 1 2 1 3079
0 7518 1 2 1 3081
0 7521 1 2 1 3125
0 7524 1 2 1 3112
0 7527 1 2 1 3063
0 7530 1 2 1 3098
0 7533 1 2 1 3133
0 7536 1 2 1 3138
0 7539 1 2 1 3150
0 7542 1 2 1 3151
0 7545 1 2 1 3162
0 7548 1 2 1 3163
0 7551 5 1 1 3338
0 7552 5 1 1 3341
0 7553 1 2 1 3230
0 7556 5 1 1 3356
0 7557 5 1 1 3358
0 7558 5 1 1 3351
0 7559 5 1 1 3353
0 7560 6 2 2 6731 6732
0 7563 6 2 2 6729 6730
0 7566 6 2 2 6735 6736
0 7569 6 2 2 6733 6734
0 7572 5 1 1 3346
0 7573 5 1 1 3348
0 7574 6 2 2 6743 6744
0 7577 6 2 2 6741 6742
0 7580 5 1 1 3360
0 7581 5 1 1 3377
0 7582 6 2 2 6753 6754
0 7585 6 2 2 6751 6752
0 7588 6 2 2 6757 6758
0 7591 6 2 2 6755 6756
0 7609 3 3 5 3096 6766 6767 6768 6769
0 7613 3 2 2 1580 6782
0 7620 3 2 5 3136 6787 6788 6789 6790
0 7649 3 1 4 3168 6836 6837 6838
0 7650 3 2 2 1622 6844
0 7655 3 3 5 3184 6848 6849 6850 6851
0 7659 3 2 2 1641 6864
0 7668 3 1 4 3210 6870 6871 6872
0 7671 3 2 5 3228 6884 6885 6886 6887
0 7744 6 1 2 2135 6968
0 7822 6 1 2 2137 7056
0 7825 3 1 4 3361 7060 7061 7062
0 7826 3 1 5 3365 7064 7065 7066 7067
0 7852 3 2 5 3370 7103 7104 7105 7106
0 8114 3 2 4 1573 6777 6778 6779
0 8117 3 2 5 1568 6770 6771 6772 6773
0 8131 4 2 3 1574 6780 6781
0 8134 4 2 4 1569 6774 6775 6776
0 8144 6 1 2 3330 7477
0 8145 6 1 2 3327 7478
0 8146 3 2 4 1617 6839 6840 6841
0 8156 4 2 3 1618 6842 6843
0 8166 3 2 4 1634 6859 6860 6861
0 8169 3 2 5 1629 6852 6853 6854 6855
0 8183 4 2 3 1635 6862 6863
0 8186 4 2 4 1630 6856 6857 6858
0 8196 3 2 4 1651 6873 6874 6875
0 8200 4 2 3 1652 6876 6877
0 8204 3 2 3 1656 6878 6879
0 8208 4 2 2 1657 6880
0 8216 6 1 2 3359 7556
0 8217 6 1 2 3357 7557
0 8218 6 1 2 3354 7558
0 8219 6 1 2 3352 7559
0 8232 6 1 2 3378 7580
0 8233 6 1 2 3376 7581
0 8242 5 1 1 4002
0 8243 5 1 1 4004
0 8244 5 1 1 4006
0 8245 5 1 1 4008
0 8246 5 1 1 4010
0 8247 5 1 1 4012
0 8248 5 1 1 4014
0 8249 5 1 1 4016
0 8250 5 1 1 4018
0 8251 5 1 1 4020
0 8252 5 1 1 3716
0 8253 5 1 1 3464
0 8254 5 1 1 3382
0 8260 5 1 1 4034
0 8261 5 1 1 4036
0 8262 7 4 2 1589 3383
0 8269 7 4 2 1611 3386
0 8274 5 1 1 3402
0 8275 5 1 1 3405
0 8276 5 1 1 3407
0 8277 5 1 1 3409
0 8278 5 1 1 3412
0 8279 5 1 1 3414
0 8280 7 1 3 2985 2982 3403
0 8281 7 1 3 3391 3388 3406
0 8282 7 1 3 2994 2991 3408
0 8283 7 1 3 3395 3393 3411
0 8284 7 1 3 3002 2999 3413
0 8285 7 1 3 3400 3397 3415
0 8288 5 1 1 3419
0 8294 5 1 1 4052
0 8295 5 1 1 4060
0 8296 5 1 1 4070
0 8297 5 1 1 4072
0 8298 7 6 2 3417 3421
0 8307 7 6 2 3422 3425
0 8315 5 1 1 4082
0 8317 5 1 1 4084
0 8319 5 1 1 4086
0 8321 5 1 1 4088
0 8322 6 1 2 4090 4543
0 8323 5 1 1 4091
0 8324 6 1 2 4092 5943
0 8325 5 1 1 4093
0 8326 6 6 2 6967 7744
0 8333 7 3 4 3435 3465 3449 3427
0 8337 7 1 2 3429 2413
0 8338 7 1 3 3437 3430 2416
0 8339 7 1 4 3450 3431 2444 3438
0 8340 7 1 2 3439 2417
0 8341 7 1 3 3451 2445 3441
0 8342 7 1 3 3467 3455 3442
0 8343 7 1 2 3443 2438
0 8344 7 1 3 2447 3456 3445
0 8345 7 1 2 3457 2448
0 8346 7 1 2 3468 3459
0 8347 7 1 2 3460 2449
0 8348 7 1 2 3471 2451
0 8349 7 1 3 3479 3472 2453
0 8350 7 1 4 3492 3473 2457 3480
0 8351 7 1 5 3506 3494 3475 3223 3481
0 8352 7 1 2 3483 2455
0 8353 7 1 3 3495 2459 3484
0 8354 7 1 4 3508 3497 3224 3485
0 8355 7 1 2 2460 3498
0 8356 7 1 3 3509 3500 3225
0 8357 7 1 2 3511 3226
0 8358 6 6 2 7055 7822
0 8365 7 3 4 3629 3541 3528 3519
0 8369 7 1 2 3520 2463
0 8370 7 1 3 3529 3522 2467
0 8371 7 1 4 3543 3523 2473 3531
0 8372 7 1 2 3532 2468
0 8373 7 1 3 3544 2475 3533
0 8374 7 1 3 3630 3546 3534
0 8375 7 1 2 3536 2469
0 8376 7 1 3 3547 2476 3537
0 8377 7 1 2 3549 2477
0 8378 7 1 2 3556 2479
0 8379 7 1 3 3567 3558 2483
0 8380 7 1 4 3588 3559 2489 3568
0 8381 7 1 5 3611 3590 3561 3231 3572
0 8382 7 1 2 3573 2484
0 8383 7 1 3 3591 2490 3575
0 8384 7 1 4 3612 3593 3233 3576
0 8385 7 1 2 3578 2485
0 8386 7 1 3 3594 2491 3579
0 8387 7 1 4 3614 3596 3234 3581
0 8388 7 1 2 3597 2492
0 8389 7 1 3 3615 3599 3235
0 8390 7 1 2 3600 2493
0 8391 7 1 3 3617 3602 3237
0 8392 7 1 2 3618 3238
0 8393 7 1 2 3632 3550
0 8394 7 9 2 3636 7063
0 8404 7 1 2 3638 7826
0 8405 7 3 4 7098 3650 3645 3639
0 8409 7 1 2 3641 4632
0 8410 7 1 3 3647 3642 4634
0 8411 7 1 4 3651 3644 4635 3648
0 8412 7 2 5 7099 3671 3666 3660 3653
0 8415 7 1 2 3654 4638
0 8416 7 1 3 3662 3656 4639
0 8417 7 1 4 3668 3657 4640 3663
0 8418 7 1 5 3672 3669 3659 4641 3665
0 8421 7 8 2 1776 3674
0 8430 7 2 4 3686 3717 3701 3677
0 8433 7 1 2 3678 2495
0 8434 7 1 3 3687 3680 2499
0 8435 7 1 4 3702 3681 2506 3689
0 8436 7 1 2 3690 2500
0 8437 7 1 3 3704 2507 3692
0 8438 7 1 3 3719 3705 3693
0 8439 7 1 2 3695 2501
0 8440 7 1 3 2509 3707 3696
0 8441 7 1 2 3708 2510
0 8442 7 1 2 3720 3710
0 8443 7 1 2 3711 2511
0 8444 7 2 5 3732 3774 3746 3723 3761
0 8447 7 1 2 3725 2512
0 8448 7 1 3 3734 3726 2514
0 8449 7 1 4 3747 3728 2517 3735
0 8450 7 1 5 3762 3749 3729 2521 3737
0 8451 7 1 2 3738 2515
0 8452 7 1 3 3750 2518 3740
0 8453 7 1 4 3764 3752 2522 3741
0 8454 7 1 2 2519 3753
0 8455 7 1 3 3765 3755 2524
0 8456 7 1 2 3767 2525
0 8457 5 2 1 3791
0 8460 5 2 1 3796
0 8463 5 2 1 3803
0 8466 5 2 1 3808
0 8469 5 1 1 3815
0 8470 5 1 1 3818
0 8471 1 2 1 3800
0 8474 1 2 1 3802
0 8477 1 2 1 3812
0 8480 1 2 1 3814
0 8483 7 1 3 3290 3286 3817
0 8484 7 1 3 3788 3785 3820
0 8485 7 2 4 3917 3845 3830 3821
0 8488 7 1 2 3823 2527
0 8489 7 1 3 3832 3824 2530
0 8490 7 1 4 3847 3826 2536 3833
0 8491 7 1 2 3835 2531
0 8492 7 1 3 3848 2539 3836
0 8493 7 1 3 3918 3850 3838
0 8494 7 1 2 3839 2532
0 8495 7 1 3 3851 2540 3841
0 8496 7 1 2 3853 2541
0 8497 7 2 5 3922 3905 3889 3869 3859
0 8500 7 1 2 3860 2543
0 8501 7 1 3 3871 3862 2547
0 8502 7 1 4 3890 3863 2553 3872
0 8503 7 1 5 3906 3892 3865 2562 3874
0 8504 7 1 2 3875 2548
0 8505 7 1 3 3893 2555 3877
0 8506 7 1 4 3907 3894 2563 3878
0 8507 7 1 4 3923 3895 3880 3908
0 8508 7 1 2 3881 2549
0 8509 7 1 3 3896 2556 3883
0 8510 7 1 4 3909 3897 2564 3884
0 8511 7 1 2 3898 2557
0 8512 7 1 3 3910 3899 2565
0 8513 7 1 3 3924 3900 3911
0 8514 7 1 2 3901 2558
0 8515 7 1 3 3912 3902 2566
0 8516 7 1 2 3913 2568
0 8517 7 1 2 3919 3854
0 8518 7 1 2 3925 3914
0 8519 5 2 1 3928
0 8522 5 2 1 3931
0 8525 1 2 1 3934
0 8528 1 2 1 3935
0 8531 1 2 1 3940
0 8534 1 2 1 3941
0 8537 5 1 1 3946
0 8538 5 1 1 3948
0 8539 7 1 3 3308 3304 3947
0 8540 7 1 3 3944 3942 3949
0 8541 7 3 4 7376 3962 3959 3950
0 8545 7 1 2 3951 4757
0 8546 7 1 3 3960 3952 4758
0 8547 7 1 4 3963 3957 4759 3961
0 8548 7 2 5 7377 3977 3974 3970 3965
0 8551 7 1 2 3966 4762
0 8552 7 1 3 3971 3967 4764
0 8553 7 1 4 3975 3968 4766 3972
0 8554 7 1 5 3978 3976 3969 4767 3973
0 8555 5 2 1 3985
0 8558 5 2 1 3990
0 8561 5 2 1 3993
0 8564 5 1 1 3998
0 8565 5 1 1 4000
0 8566 1 2 1 3988
0 8569 1 2 1 3989
0 8572 1 2 1 3996
0 8575 1 2 1 3997
0 8578 7 1 3 3318 3314 3999
0 8579 7 1 3 3981 3979 4001
0 8580 1 2 1 3776
0 8583 1 2 1 3731
0 8586 1 2 1 3743
0 8589 1 2 1 3756
0 8592 1 2 1 3768
0 8595 1 2 1 3476
0 8598 1 2 1 3488
0 8601 1 2 1 3501
0 8604 1 2 1 3512
0 8607 5 1 1 4022
0 8608 6 1 2 4023 5469
0 8609 5 1 1 4024
0 8610 6 1 2 4025 4793
0 8615 5 1 1 4026
0 8616 5 1 1 4028
0 8617 5 1 1 4030
0 8618 5 1 1 4032
0 8619 5 1 1 4044
0 8624 5 1 1 4038
0 8625 5 1 1 4040
0 8626 5 1 1 4042
0 8627 6 2 2 8144 8145
0 8632 5 1 1 4046
0 8633 5 1 1 4048
0 8634 5 1 1 4050
0 8637 5 1 1 4054
0 8638 5 1 1 4056
0 8639 5 1 1 4058
0 8644 5 1 1 4062
0 8645 5 1 1 4064
0 8646 5 1 1 4066
0 8647 5 1 1 4068
0 8648 5 1 1 4080
0 8653 5 1 1 4074
0 8654 5 1 1 4076
0 8655 5 1 1 4078
0 8660 1 2 1 3433
0 8663 1 2 1 3434
0 8666 1 2 1 3446
0 8669 1 2 1 3447
0 8672 1 2 1 3461
0 8675 1 2 1 3463
0 8678 1 2 1 3633
0 8681 1 2 1 3554
0 8684 1 2 1 3525
0 8687 1 2 1 3538
0 8690 1 2 1 3635
0 8693 1 2 1 3555
0 8696 1 2 1 3526
0 8699 1 2 1 3540
0 8702 1 2 1 3620
0 8705 1 2 1 3562
0 8708 1 2 1 3603
0 8711 1 2 1 3582
0 8714 1 2 1 3584
0 8717 5 1 1 4094
0 8718 1 2 1 3621
0 8721 1 2 1 3564
0 8724 1 2 1 3605
0 8727 6 2 2 8216 8217
0 8730 6 2 2 8218 8219
0 8733 5 1 1 4104
0 8734 5 1 1 4106
0 8735 1 2 1 3683
0 8738 1 2 1 3684
0 8741 1 2 1 3698
0 8744 1 2 1 3699
0 8747 1 2 1 3713
0 8750 1 2 1 3714
0 8753 5 1 1 4096
0 8754 5 1 1 4098
0 8755 5 1 1 4100
0 8756 5 1 1 4102
0 8757 1 2 1 3920
0 8760 1 2 1 3856
0 8763 1 2 1 3827
0 8766 1 2 1 3842
0 8769 1 2 1 3921
0 8772 1 2 1 3857
0 8775 1 2 1 3829
0 8778 1 2 1 3844
0 8781 1 2 1 3926
0 8784 1 2 1 3915
0 8787 1 2 1 3866
0 8790 1 2 1 3903
0 8793 1 2 1 3886
0 8796 1 2 1 3887
0 8799 1 2 1 3927
0 8802 1 2 1 3916
0 8805 1 2 1 3868
0 8808 1 2 1 3904
0 8811 6 2 2 8232 8233
0 8814 5 1 1 4112
0 8815 5 1 1 4114
0 8816 5 1 1 4108
0 8817 5 1 1 4110
0 8818 7 1 2 4121 1612
0 8840 7 1 2 1590 4116
0 8857 5 3 1 4117
0 8861 7 1 3 3389 2986 8274
0 8862 7 1 3 2983 3392 8275
0 8863 7 1 3 3394 2995 8276
0 8864 7 1 3 2992 3396 8277
0 8865 7 1 3 3399 3003 8278
0 8866 7 1 3 3000 3401 8279
0 8871 5 2 1 4125
0 8874 7 1 2 3418 4126
0 8878 7 1 2 4130 3423
0 8879 5 1 1 4154
0 8880 6 1 2 4155 8315
0 8881 5 1 1 4156
0 8882 6 1 2 4157 8317
0 8883 5 1 1 4158
0 8884 6 1 2 4159 8319
0 8885 5 1 1 4160
0 8886 6 1 2 4161 8321
0 8887 6 1 2 2133 8323
0 8888 6 1 2 2590 8325
0 8898 3 3 4 4544 8337 8338 8339
0 8902 3 2 5 4562 8348 8349 8350 8351
0 8920 3 3 4 4576 8369 8370 8371
0 8924 3 2 2 2471 8377
0 8927 3 3 5 4592 8378 8379 8380 8381
0 8931 3 2 2 2494 8392
0 8943 3 3 2 7825 8404
0 8950 3 3 4 4630 8409 8410 8411
0 8956 3 2 5 4637 8415 8416 8417 8418
0 8959 5 1 1 4132
0 8960 7 1 2 1777 4133
0 8963 3 1 4 4656 8433 8434 8435
0 8966 3 2 5 4674 8447 8448 8449 8450
0 8991 7 1 3 3787 3291 8469
0 8992 7 1 3 3288 3790 8470
0 8995 3 1 4 4701 8488 8489 8490
0 8996 3 2 2 2534 8496
0 9001 3 3 5 4717 8500 8501 8502 8503
0 9005 3 2 2 2559 8516
0 9024 7 1 3 3943 3309 8537
0 9025 7 1 3 3305 3945 8538
0 9029 3 3 4 4756 8545 8546 8547
0 9035 3 2 5 4760 8551 8552 8553 8554
0 9053 7 1 3 3980 3319 8564
0 9054 7 1 3 3316 3982 8565
0 9064 6 1 2 2411 8607
0 9065 6 1 2 1987 8609
0 9066 5 1 1 4134
0 9067 6 1 2 4135 4795
0 9068 3 2 2 4119 6783
0 9071 5 1 1 4136
0 9072 5 1 1 4138
0 9073 6 1 2 4139 6195
0 9074 5 2 1 4120
0 9077 5 1 1 4140
0 9079 3 2 2 4123 6865
0 9082 5 1 1 4142
0 9083 5 2 1 4124
0 9086 5 1 1 4144
0 9087 5 1 1 4146
0 9088 6 1 2 4147 4813
0 9089 3 2 2 4128 6866
0 9092 5 1 1 4148
0 9093 5 1 1 4150
0 9094 6 1 2 4151 6203
0 9095 5 2 1 4129
0 9098 5 1 1 4152
0 9099 3 2 4 2414 8340 8341 8342
0 9103 4 2 3 2415 8343 8344
0 9107 3 2 3 2439 8345 8346
0 9111 4 2 2 2440 8347
0 9117 3 2 4 2464 8372 8373 8374
0 9127 4 2 3 2465 8375 8376
0 9146 4 2 3 2486 8390 8391
0 9149 4 2 4 2480 8385 8386 8387
0 9159 6 1 2 4107 8733
0 9160 6 1 2 4105 8734
0 9161 3 2 4 2497 8436 8437 8438
0 9165 4 2 3 2498 8439 8440
0 9169 3 2 3 2503 8441 8442
0 9173 4 2 2 2504 8443
0 9179 6 1 2 4099 8753
0 9180 6 1 2 4097 8754
0 9181 6 1 2 4103 8755
0 9182 6 1 2 4101 8756
0 9183 3 2 4 2528 8491 8492 8493
0 9193 4 2 3 2529 8494 8495
0 9203 3 2 4 2551 8511 8512 8513
0 9206 3 2 5 2544 8504 8505 8506 8507
0 9220 4 2 3 2552 8514 8515
0 9223 4 2 4 2545 8508 8509 8510
0 9234 6 1 2 4115 8814
0 9235 6 1 2 4113 8815
0 9236 6 1 2 4111 8816
0 9237 6 1 2 4109 8817
0 9238 3 1 2 1614 8818
0 9242 3 1 2 1592 8840
0 9243 6 1 2 8324 8888
0 9244 5 1 1 4278
0 9245 5 1 1 4280
0 9246 5 1 1 4282
0 9247 5 1 1 4284
0 9248 5 1 1 4286
0 9249 5 1 1 4288
0 9250 5 1 1 4290
0 9251 5 1 1 4292
0 9252 5 1 1 4294
0 9256 4 1 2 8861 8280
0 9257 4 1 2 8862 8281
0 9258 4 1 2 8863 8282
0 9259 4 1 2 8864 8283
0 9260 4 1 2 8865 8284
0 9261 4 1 2 8866 8285
0 9262 5 1 1 4296
0 9265 3 2 2 7649 8874
0 9268 3 2 2 7668 8878
0 9271 6 1 2 4083 8879
0 9272 6 1 2 4085 8881
0 9273 6 1 2 4087 8883
0 9274 6 1 2 4089 8885
0 9275 6 1 2 8322 8887
0 9276 5 1 1 4188
0 9280 7 2 5 3489 4182 3503 3477 3513
0 9285 7 1 5 370 4183 3504 3514 3491
0 9286 7 1 4 371 4184 3505 3516
0 9287 7 1 3 372 4185 3517
0 9288 7 1 2 373 4186
0 9290 5 1 1 4298
0 9292 5 1 1 4300
0 9294 5 1 1 4302
0 9296 5 1 1 4305
0 9297 6 1 2 4307 5966
0 9298 5 1 1 4309
0 9299 6 1 2 4310 6969
0 9300 5 1 1 4311
0 9301 5 1 1 4198
0 9307 7 3 5 4191 3623 3606 3585 3565
0 9314 7 1 4 4192 3608 3587 3624
0 9315 7 1 3 4194 3609 3626
0 9318 7 1 2 4195 3627
0 9319 5 1 1 4319
0 9320 5 1 1 4329
0 9321 5 1 1 4339
0 9322 5 1 1 4341
0 9323 5 1 1 4349
0 9324 5 1 1 4351
0 9326 5 1 1 4210
0 9332 7 6 2 4211 4213
0 9339 3 2 2 2408 8960
0 9344 7 6 2 4223 4225
0 9352 5 1 1 4353
0 9354 5 1 1 4355
0 9356 5 1 1 4357
0 9358 5 1 1 4359
0 9359 6 1 2 4361 6078
0 9360 5 1 1 4362
0 9361 6 1 2 4363 7187
0 9362 5 1 1 4364
0 9363 5 1 1 4235
0 9364 5 1 1 4237
0 9365 5 1 1 4239
0 9366 5 1 1 4241
0 9367 4 1 2 8991 8483
0 9368 4 1 2 8992 8484
0 9369 7 1 3 3797 3793 4236
0 9370 7 1 3 4229 4227 4238
0 9371 7 1 3 3809 3805 4240
0 9372 7 1 3 4233 4231 4242
0 9375 5 1 1 4245
0 9381 5 1 1 4371
0 9382 5 1 1 4379
0 9383 5 1 1 4389
0 9384 5 1 1 4391
0 9385 7 6 2 4243 4246
0 9392 5 1 1 4251
0 9393 5 1 1 4253
0 9394 5 1 1 4255
0 9395 5 1 1 4257
0 9396 7 1 3 3932 3929 4252
0 9397 7 1 3 4249 4247 4254
0 9398 7 1 3 3300 3296 4256
0 9399 7 1 3 3938 3936 4258
0 9400 4 1 2 9024 8539
0 9401 4 1 2 9025 8540
0 9402 5 1 1 4259
0 9407 6 1 2 4262 90
0 9408 7 3 2 4260 4263
0 9412 5 1 1 4401
0 9413 5 1 1 4270
0 9414 5 1 1 4272
0 9415 5 1 1 4274
0 9416 5 1 1 4276
0 9417 4 1 2 9053 8578
0 9418 4 1 2 9054 8579
0 9419 7 1 3 3986 3324 4271
0 9420 7 1 3 4264 3983 4273
0 9421 7 1 3 3994 3991 4275
0 9422 7 1 3 4268 4266 4277
0 9423 1 2 1 4187
0 9426 6 2 2 9064 8608
0 9429 6 2 2 9065 8610
0 9432 6 1 2 2000 9066
0 9435 6 1 2 2580 9072
0 9442 6 1 2 2104 9087
0 9445 6 1 2 2588 9093
0 9454 5 1 1 4312
0 9455 5 1 1 4315
0 9456 5 1 1 4317
0 9459 5 1 1 4321
0 9460 5 1 1 4323
0 9461 5 1 1 4325
0 9462 1 2 1 4196
0 9465 5 1 1 4331
0 9466 5 1 1 4335
0 9467 5 1 1 4337
0 9468 5 1 1 4347
0 9473 1 2 1 4197
0 9476 5 1 1 4343
0 9477 5 1 1 4345
0 9478 6 2 2 9159 9160
0 9485 6 2 2 9179 9180
0 9488 6 2 2 9181 9182
0 9493 5 1 1 4365
0 9494 5 1 1 4367
0 9495 5 1 1 4369
0 9498 5 1 1 4373
0 9499 5 1 1 4375
0 9500 5 1 1 4377
0 9505 5 1 1 4381
0 9506 5 1 1 4383
0 9507 5 1 1 4385
0 9508 5 1 1 4387
0 9509 5 1 1 4399
0 9514 5 1 1 4393
0 9515 5 1 1 4395
0 9516 5 1 1 4397
0 9517 6 2 2 9234 9235
0 9520 6 2 2 9236 9237
0 9526 7 1 2 4425 4215
0 9531 7 1 2 4426 4216
0 9539 6 1 2 9271 8880
0 9540 6 1 2 9273 8884
0 9541 5 1 1 9275
0 9543 7 2 2 4403 8254
0 9551 7 2 2 4406 8288
0 9555 6 1 2 9272 8882
0 9556 6 1 2 9274 8886
0 9557 5 1 1 4408
0 9560 7 1 2 4413 4189
0 9561 5 1 1 4459
0 9562 6 1 2 4460 9290
0 9563 5 1 1 4461
0 9564 6 1 2 4462 9292
0 9565 5 1 1 4546
0 9566 6 1 2 4547 9294
0 9567 5 1 1 4548
0 9568 6 1 2 4550 9296
0 9569 6 1 2 2610 9298
0 9570 6 1 2 3335 9300
0 9571 5 1 1 4415
0 9575 5 3 1 4420
0 9579 7 1 2 4199 4421
0 9581 5 1 1 4428
0 9582 5 1 1 4431
0 9585 7 1 2 4212 4432
0 9591 7 1 2 4433 4224
0 9592 5 1 1 4560
0 9593 6 1 2 4561 9352
0 9594 5 1 1 4564
0 9595 6 1 2 4565 9354
0 9596 5 1 1 4567
0 9597 6 1 2 4568 9356
0 9598 5 1 1 4569
0 9599 6 1 2 4571 9358
0 9600 6 1 2 2691 9360
0 9601 6 1 2 3345 9362
0 9602 7 1 3 4228 3799 9363
0 9603 7 1 3 3794 4230 9364
0 9604 7 1 3 4232 3811 9365
0 9605 7 1 3 3806 4234 9366
0 9608 5 2 1 4437
0 9611 7 1 2 4244 4438
0 9612 7 1 3 4248 3933 9392
0 9613 7 1 3 3930 4250 9393
0 9614 7 1 3 3937 3301 9394
0 9615 7 1 3 3297 3939 9395
0 9616 5 1 1 4442
0 9617 5 1 1 4445
0 9618 7 1 2 4261 4446
0 9621 7 1 3 3984 3987 9413
0 9622 7 1 3 3325 4265 9414
0 9623 7 1 3 4267 3995 9415
0 9624 7 1 3 3992 4269 9416
0 9626 3 2 5 2452 8352 8353 8354 9285
0 9629 3 2 4 2456 8355 8356 9286
0 9632 3 2 3 2461 8357 9287
0 9635 3 2 2 3227 9288
0 9642 6 2 2 9067 9432
0 9645 5 1 1 4447
0 9646 6 2 2 9073 9435
0 9649 5 1 1 4449
0 9650 6 2 2 9257 9256
0 9653 6 2 2 9259 9258
0 9656 6 2 2 9261 9260
0 9659 5 1 1 4451
0 9660 6 1 2 4452 4809
0 9661 5 1 1 4453
0 9662 6 1 2 4454 6202
0 9663 6 2 2 9088 9442
0 9666 5 1 1 4455
0 9667 6 2 2 9094 9445
0 9670 5 1 1 4457
0 9671 3 2 2 4418 8393
0 9674 5 1 1 4551
0 9675 5 2 1 4419
0 9678 5 1 1 4553
0 9679 3 2 4 2487 8388 8389 9315
0 9682 3 2 2 4423 9318
0 9685 3 2 5 2481 8382 8383 8384 9314
0 9690 5 1 1 4556
0 9691 6 1 2 4557 8717
0 9692 5 2 1 4424
0 9695 5 1 1 4558
0 9698 6 2 2 9401 9400
0 9702 6 2 2 9368 9367
0 9707 3 2 2 4435 8517
0 9710 5 1 1 4572
0 9711 5 2 1 4436
0 9714 5 1 1 4574
0 9715 5 1 1 4579
0 9716 6 1 2 4580 6235
0 9717 3 2 2 4440 8518
0 9720 5 1 1 4582
0 9721 5 1 1 4584
0 9722 6 1 2 4585 7573
0 9723 5 2 1 4441
0 9726 5 1 1 4587
0 9727 6 2 2 9418 9417
0 9732 7 1 2 4591 4166
0 9733 6 1 2 9581 9326
0 9734 7 1 5 91 4670 4601 4201 4217
0 9735 7 1 5 92 4671 4602 4202 4218
0 9736 7 1 2 4589 4162
0 9737 5 1 1 9555
0 9738 5 1 1 9556
0 9739 6 1 2 9361 9601
0 9740 6 1 2 4673 1115
0 9741 5 1 1 4676
0 9742 6 1 2 9299 9570
0 9754 7 3 2 4190 4595
0 9758 3 3 2 4409 9560
0 9762 6 1 2 4299 9561
0 9763 6 1 2 4301 9563
0 9764 6 1 2 4304 9565
0 9765 6 1 2 4306 9567
0 9766 6 1 2 9297 9569
0 9767 7 1 2 4596 374
0 9768 6 1 2 9557 9276
0 9769 5 1 1 4598
0 9773 6 1 2 4599 375
0 9774 6 1 2 9571 9301
0 9775 7 3 2 4200 4600
0 9779 3 3 2 4416 9579
0 9784 5 1 1 4688
0 9785 6 1 2 9616 9402
0 9786 3 3 2 4429 9585
0 9790 7 1 4 93 4672 4604 4203
0 9791 3 3 2 8963 9591
0 9795 6 1 2 4354 9592
0 9796 6 1 2 4356 9594
0 9797 6 1 2 4358 9596
0 9798 6 1 2 4360 9598
0 9799 6 1 2 9359 9600
0 9800 4 1 2 9602 9369
0 9801 4 1 2 9603 9370
0 9802 4 1 2 9604 9371
0 9803 4 1 2 9605 9372
0 9805 5 1 1 4690
0 9806 5 1 1 4692
0 9809 3 3 2 8995 9611
0 9813 4 1 2 9612 9396
0 9814 4 1 2 9613 9397
0 9815 4 1 2 9614 9398
0 9816 4 1 2 9615 9399
0 9817 7 2 2 9617 9407
0 9820 3 3 2 4443 9618
0 9825 5 1 1 4704
0 9826 5 1 1 4707
0 9827 4 1 2 9621 9419
0 9828 4 1 2 9622 9420
0 9829 4 1 2 9623 9421
0 9830 4 1 2 9624 9422
0 9835 5 1 1 4677
0 9836 6 1 2 4679 4789
0 9837 5 1 1 4680
0 9838 6 1 2 4681 4794
0 9846 6 1 2 2102 9659
0 9847 6 1 2 2586 9661
0 9862 5 1 1 4683
0 9863 6 1 2 4095 9690
0 9866 5 1 1 4685
0 9873 6 1 2 2767 9715
0 9876 6 1 2 3350 9721
0 9890 6 1 2 9795 9593
0 9891 6 1 2 9797 9597
0 9892 5 1 1 9799
0 9893 6 1 2 680 9741
0 9894 6 1 2 9762 9562
0 9895 6 1 2 9764 9566
0 9896 5 1 1 9766
0 9897 5 1 1 4721
0 9898 6 1 2 4723 9249
0 9899 5 1 1 4724
0 9900 6 1 2 4725 9250
0 9901 5 1 1 4726
0 9902 6 1 2 4727 9251
0 9903 5 1 1 4729
0 9904 6 1 2 4730 9252
0 9905 5 1 1 4709
0 9906 5 1 1 4736
0 9907 6 1 2 4737 5769
0 9908 5 1 1 4738
0 9909 6 1 2 4739 5770
0 9910 5 1 1 4740
0 9911 6 1 2 4741 9262
0 9917 5 1 1 4712
0 9923 6 1 2 9763 9564
0 9924 6 1 2 9765 9568
0 9925 3 6 2 4414 9767
0 9932 7 2 2 4714 9773
0 9935 7 2 2 4715 9769
0 9938 5 1 1 4807
0 9939 6 1 2 4808 9323
0 9945 6 1 2 9796 9595
0 9946 6 1 2 9798 9599
0 9947 5 1 1 4811
0 9948 6 1 2 4812 6102
0 9949 7 2 2 4719 9375
0 9953 5 1 1 4827
0 9954 6 1 2 4828 9412
0 9955 6 1 2 1985 9835
0 9956 6 1 2 1998 9837
0 9957 5 1 1 4731
0 9958 6 1 2 4732 9645
0 9959 5 1 1 4733
0 9960 6 1 2 4734 9649
0 9961 6 2 2 9660 9846
0 9964 6 2 2 9662 9847
0 9967 5 1 1 4742
0 9968 6 1 2 4770 9666
0 9969 5 1 1 4771
0 9970 6 1 2 4772 9670
0 9971 5 1 1 4773
0 9972 6 1 2 4774 6213
0 9973 5 1 1 4785
0 9974 6 1 2 4786 7551
0 9975 5 1 1 4787
0 9976 6 1 2 4788 7552
0 9977 5 1 1 4791
0 9978 5 1 1 4797
0 9979 6 2 2 9691 9863
0 9982 5 1 1 4804
0 9983 6 2 2 9814 9813
0 9986 6 2 2 9816 9815
0 9989 6 2 2 9801 9800
0 9992 6 2 2 9803 9802
0 9995 5 1 1 4815
0 9996 6 1 2 4816 6231
0 9997 5 1 1 4818
0 9998 6 1 2 4819 7572
0 9999 6 2 2 9716 9873
0 10002 5 1 1 4821
0 10003 6 2 2 9722 9876
0 10006 5 1 1 4824
0 10007 6 2 2 9830 9829
0 10010 6 2 2 9828 9827
0 10013 7 1 3 4852 4176 4167
0 10014 7 1 4 4834 4654 4177 4168
0 10015 7 1 5 376 4830 4655 4178 4169
0 10016 7 1 3 4848 4204 4219
0 10017 7 1 4 4864 4605 4205 4220
0 10018 7 1 3 4849 4206 4221
0 10019 7 1 4 4866 4606 4207 4222
0 10020 7 1 3 4857 4170 4163
0 10021 7 1 4 4843 4663 4171 4164
0 10022 7 1 5 377 4839 4664 4172 4165
0 10023 5 1 1 9945
0 10024 5 1 1 9946
3 10025 6 0 2 9740 9893
0 10026 5 1 1 9923
0 10028 5 1 1 9924
0 10032 6 1 2 4289 9897
0 10033 6 1 2 4291 9899
0 10034 6 1 2 4293 9901
0 10035 6 1 2 4295 9903
0 10036 6 1 2 2582 9906
0 10037 6 1 2 2584 9908
0 10038 6 1 2 4297 9910
0 10039 7 1 2 4858 4173
0 10040 7 1 3 4845 4665 4174
0 10041 7 1 4 378 4840 4666 4175
0 10042 7 1 2 4846 4668
0 10043 7 1 3 379 4842 4669
0 10050 6 1 2 4350 9938
0 10053 5 1 1 4861
0 10054 7 1 2 4863 4444
0 10055 7 1 2 4851 4208
0 10056 7 1 3 4867 4607 4209
0 10057 7 1 2 4854 4179
0 10058 7 1 3 4836 4658 4180
0 10059 7 1 4 380 4831 4659 4181
0 10060 7 1 2 4837 4660
0 10061 7 1 3 381 4833 4662
0 10062 6 1 2 2736 9947
0 10067 6 1 2 4402 9953
0 10070 6 2 2 9955 9836
0 10073 6 2 2 9956 9838
0 10076 6 1 2 4448 9957
0 10077 6 1 2 4450 9959
0 10082 6 1 2 4456 9967
0 10083 6 1 2 4458 9969
0 10084 6 1 2 2633 9971
0 10085 6 1 2 3339 9973
0 10086 6 1 2 3342 9975
0 10093 6 1 2 2763 9995
0 10094 6 1 2 3347 9997
3 10101 3 0 5 9238 9732 10013 10014 10015
3 10102 3 0 5 4608 9526 10016 10017 9734
3 10103 3 0 5 4609 9531 10018 10019 9735
3 10104 3 0 5 9242 9736 10020 10021 10022
0 10105 7 1 2 4869 9894
0 10106 7 1 2 4870 9895
0 10107 7 1 2 4872 9896
0 10108 7 1 2 4873 8253
3 10109 6 0 2 10032 9898
3 10110 6 0 2 10033 9900
3 10111 6 0 2 10034 9902
3 10112 6 0 2 10035 9904
0 10113 6 1 2 10036 9907
0 10114 6 1 2 10037 9909
0 10115 6 1 2 10038 9911
0 10116 3 2 4 4590 10039 10040 10041
0 10119 3 4 3 4860 10042 10043
0 10124 5 5 1 4875
0 10130 7 1 2 9768 4876
0 10131 5 1 1 4878
0 10132 5 1 1 4881
0 10133 7 1 2 4879 4417
0 10134 6 1 2 10050 9939
0 10135 5 1 1 4896
0 10136 6 1 2 4897 9324
0 10137 5 1 1 4899
0 10138 6 1 2 4900 9784
0 10139 7 1 2 9785 10053
0 10140 3 1 4 4427 10055 10056 9790
0 10141 3 6 4 4594 10057 10058 10059
0 10148 3 6 3 4855 10060 10061
0 10155 6 1 2 10062 9948
0 10156 5 1 1 4902
0 10157 6 1 2 4903 9805
0 10158 5 1 1 4905
0 10159 6 1 2 4906 9806
0 10160 5 1 1 4884
0 10161 6 1 2 10067 9954
0 10162 5 1 1 4914
0 10163 6 1 2 4915 9825
0 10164 5 1 1 4917
0 10165 6 1 2 4918 9826
0 10170 6 2 2 10076 9958
0 10173 6 2 2 10077 9960
0 10176 5 1 1 4887
0 10177 6 1 2 4888 9082
0 10178 5 1 1 4890
0 10179 6 1 2 4891 9086
0 10180 6 2 2 10082 9968
0 10183 6 2 2 10083 9970
0 10186 6 2 2 9972 10084
0 10189 6 2 2 9974 10085
0 10192 6 2 2 9976 10086
0 10195 5 1 1 4893
0 10196 6 1 2 4894 9982
0 10197 6 2 2 9996 10093
0 10200 6 2 2 9998 10094
0 10203 5 1 1 4908
0 10204 6 1 2 4909 10002
0 10205 5 1 1 4911
0 10206 6 1 2 4912 10006
0 10212 6 1 2 4920 4308
0 10213 6 1 2 4923 4313
0 10230 7 1 2 9774 10131
0 10231 6 1 2 4352 10135
0 10232 6 1 2 4689 10137
0 10233 3 1 2 10139 10054
0 10234 6 1 2 3675 10140
0 10237 6 1 2 4691 10156
0 10238 6 1 2 4703 10158
0 10239 6 1 2 4705 10162
0 10240 6 1 2 4708 10164
0 10241 5 1 1 4921
0 10242 5 1 1 4924
0 10247 6 1 2 4143 10176
0 10248 6 1 2 4145 10178
0 10259 6 1 2 4805 10195
0 10264 6 1 2 4822 10203
0 10265 6 1 2 4825 10205
0 10266 7 1 2 10026 4935
0 10267 7 1 2 10028 4936
0 10268 7 1 2 9742 4938
0 10269 7 1 2 3469 4939
0 10270 6 1 2 3385 4926
0 10271 6 1 2 1556 10241
0 10272 6 1 2 1558 10242
0 10273 1 4 1 4927
0 10278 7 1 5 4942 2977 2964 2972 2955
0 10279 7 1 4 4944 2978 2965 2973
0 10280 7 1 3 4945 2979 2974
0 10281 7 1 2 4947 2980
0 10282 7 1 2 3387 4948
0 10283 5 3 1 4929
0 10287 7 1 5 4951 3218 3201 3212 3191
0 10288 7 1 4 4953 3219 3203 3213
0 10289 7 1 3 4954 3220 3214
0 10290 7 1 2 4956 3222
0 10291 7 1 2 3426 4957
0 10292 7 1 2 4410 4941
0 10293 6 1 2 10231 10136
0 10294 6 1 2 10232 10138
0 10295 6 1 2 4214 10233
0 10296 7 2 2 8959 10234
0 10299 6 1 2 10237 10157
0 10300 6 1 2 10238 10159
0 10301 3 4 2 10230 10133
0 10306 6 1 2 10239 10163
0 10307 6 1 2 10240 10165
0 10308 1 2 1 4959
0 10311 1 2 1 4950
0 10314 5 1 1 4960
0 10315 6 1 2 4962 9071
0 10316 5 1 1 4963
0 10317 6 1 2 4965 9077
0 10318 6 2 2 10247 10177
0 10321 6 2 2 10248 10179
0 10324 5 1 1 4966
0 10325 6 1 2 4968 9092
0 10326 5 1 1 4969
0 10327 6 1 2 4971 9098
0 10328 5 1 1 4972
0 10329 6 1 2 4974 9674
0 10330 5 1 1 4975
0 10331 6 1 2 4977 9678
0 10332 5 1 1 4978
0 10333 6 1 2 4980 9977
0 10334 6 2 2 10259 10196
0 10337 5 1 1 4981
0 10338 6 1 2 4983 9710
0 10339 5 1 1 4984
0 10340 6 1 2 4986 9714
0 10341 6 2 2 10264 10204
0 10344 6 2 2 10265 10206
3 10350 3 0 2 10266 10105
3 10351 3 0 2 10267 10106
3 10352 3 0 2 10268 10107
3 10353 3 0 2 10269 10108
0 10354 7 2 2 4404 10270
0 10357 6 2 2 10271 10212
0 10360 6 2 2 10272 10213
0 10367 3 4 2 4122 10282
0 10375 3 5 2 4131 10291
0 10381 3 6 2 10292 10130
0 10388 7 2 4 10114 10134 10293 10294
0 10391 7 2 2 9582 10295
0 10399 7 2 4 10113 10115 10299 10300
0 10402 7 2 4 10155 10161 10306 10307
0 10406 3 2 5 1665 6888 6889 6890 10287
0 10409 3 2 4 1668 6891 6892 10288
0 10412 3 2 3 1672 6893 10289
0 10415 3 2 2 1677 10290
0 10419 3 2 5 1597 6791 6792 6793 10278
0 10422 3 2 4 1600 6794 6795 10279
0 10425 3 2 3 1604 6796 10280
0 10428 3 2 2 1609 10281
0 10431 6 1 2 4137 10314
0 10432 6 1 2 4141 10316
0 10437 6 1 2 4149 10324
0 10438 6 1 2 4153 10326
0 10439 6 1 2 4552 10328
0 10440 6 1 2 4554 10330
0 10441 6 1 2 4792 10332
0 10444 6 1 2 4573 10337
0 10445 6 1 2 4578 10339
0 10450 5 1 1 4998
0 10451 7 1 2 4999 2409
0 10455 5 1 1 5007
0 10456 6 1 2 5008 8242
0 10465 5 1 1 5010
0 10466 6 1 2 5011 8247
0 10479 5 3 1 4987
0 10497 5 3 1 5001
0 10509 6 2 2 10431 10315
0 10512 6 2 2 10432 10317
0 10515 5 1 1 5013
0 10516 6 1 2 5014 8632
0 10517 5 1 1 5016
0 10518 6 1 2 5017 8637
0 10519 6 2 2 10437 10325
0 10522 6 2 2 10438 10327
0 10525 6 2 2 10439 10329
0 10528 6 2 2 10440 10331
0 10531 6 2 2 10441 10333
0 10534 5 1 1 5019
0 10535 6 1 2 5020 9695
0 10536 6 2 2 10444 10338
0 10539 6 2 2 10445 10340
0 10542 5 1 1 5022
0 10543 6 1 2 5023 9720
0 10544 5 1 1 5025
0 10545 6 1 2 5026 9726
0 10546 7 1 2 5631 10450
0 10547 5 1 1 5070
0 10548 7 1 2 5072 4430
0 10549 7 1 2 5165 5037
0 10550 5 1 1 5028
0 10551 7 1 2 5029 1593
0 10552 6 1 2 4003 10455
0 10553 7 1 2 5043 9539
0 10554 7 1 2 5044 9540
0 10555 7 1 2 5050 9541
0 10556 7 1 2 5051 6761
0 10557 5 1 1 5079
0 10558 6 1 2 5081 8243
0 10559 5 1 1 5082
0 10560 6 1 2 5084 8244
0 10561 5 1 1 5085
0 10562 6 1 2 5087 8245
0 10563 5 1 1 5088
0 10564 6 1 2 5090 8246
0 10565 6 1 2 4013 10465
0 10566 5 1 1 5091
0 10567 6 1 2 5093 8248
0 10568 5 1 1 5094
0 10569 6 1 2 5096 8249
0 10570 5 1 1 5097
0 10571 6 1 2 5099 8250
0 10572 5 1 1 5100
0 10573 6 1 2 5102 8251
3 10574 5 0 1 5073
3 10575 5 0 1 5076
3 10576 5 0 1 5063
0 10577 7 1 3 5075 5078 5069
0 10581 7 1 3 5034 4710 4989
0 10582 7 1 3 5031 9905 4990
0 10583 5 3 1 5038
0 10587 7 1 2 5040 5735
0 10588 7 1 2 5041 3135
0 10589 5 4 1 5053
0 10594 7 1 5 5054 3777 3758 3770 3744
0 10595 7 1 4 5056 3779 3759 3771
0 10596 7 1 3 5057 3780 3773
0 10597 7 1 2 5059 3784
0 10598 7 1 2 4226 5060
0 10602 1 2 1 5062
0 10609 6 1 2 4047 10515
0 10610 6 1 2 4055 10517
0 10621 6 1 2 4559 10534
0 10626 6 1 2 4583 10542
0 10627 6 1 2 4588 10544
3 10628 3 0 2 10546 10451
0 10629 7 1 2 9733 10547
0 10631 7 1 2 5166 10550
3 10632 6 0 2 10552 10456
0 10637 6 1 2 4005 10557
0 10638 6 1 2 4007 10559
0 10639 6 1 2 4009 10561
0 10640 6 1 2 4011 10563
3 10641 6 0 2 10565 10466
0 10642 6 1 2 4015 10566
0 10643 6 1 2 4017 10568
0 10644 6 1 2 4019 10570
0 10645 6 1 2 4021 10572
0 10647 7 1 3 886 887 10577
0 10648 7 1 3 5035 4405 5103
0 10649 7 1 3 5032 4118 5105
0 10652 3 5 2 4434 10598
0 10659 3 2 5 2513 8451 8452 8453 10594
0 10662 3 2 4 2516 8454 8455 10595
0 10665 3 2 3 2520 8456 10596
0 10668 3 2 2 2526 10597
0 10671 5 1 1 5116
0 10672 6 1 2 5118 8615
0 10673 5 1 1 5119
0 10674 6 1 2 5121 8624
0 10675 6 2 2 10609 10516
0 10678 6 2 2 10610 10518
0 10681 5 1 1 5122
0 10682 6 1 2 5124 8644
0 10683 5 1 1 5125
0 10684 6 1 2 5127 8653
0 10685 5 1 1 5128
0 10686 6 1 2 5130 9454
0 10687 5 1 1 5131
0 10688 6 1 2 5133 9459
0 10689 5 1 1 5134
0 10690 6 1 2 5136 9978
0 10691 6 2 2 10621 10535
0 10694 5 1 1 5137
0 10695 6 1 2 5139 9493
0 10696 5 1 1 5140
0 10697 6 1 2 5142 9498
0 10698 6 2 2 10626 10543
0 10701 6 2 2 10627 10545
3 10704 3 0 2 10629 10548
0 10705 7 1 2 1615 5143
3 10706 3 0 2 10631 10551
0 10707 7 1 2 9737 5148
0 10708 7 1 2 9738 5149
0 10709 7 1 2 9243 5151
0 10710 7 1 2 3171 5152
3 10711 6 0 2 10637 10558
3 10712 6 0 2 10638 10560
3 10713 6 0 2 10639 10562
3 10714 6 0 2 10640 10564
3 10715 6 0 2 10642 10567
3 10716 6 0 2 10643 10569
3 10717 6 0 2 10644 10571
3 10718 6 0 2 10645 10573
0 10719 5 1 1 5154
0 10720 6 1 2 5155 9244
3 10729 5 0 1 10647
0 10730 7 1 2 5178 5145
0 10731 7 1 2 1345 5146
0 10737 6 1 2 4027 10671
0 10738 6 1 2 4039 10673
0 10739 3 2 4 10648 10649 10581 10582
0 10746 6 1 2 4063 10681
0 10747 6 1 2 4075 10683
0 10748 6 1 2 4314 10685
0 10749 6 1 2 4322 10687
0 10750 6 1 2 4798 10689
0 10753 6 1 2 4366 10694
0 10754 6 1 2 4374 10696
3 10759 3 0 2 10705 10549
3 10760 3 0 2 10707 10553
3 10761 3 0 2 10708 10554
3 10762 3 0 2 10709 10555
3 10763 3 0 2 10710 10556
0 10764 6 1 2 4279 10719
0 10765 7 1 2 5157 9890
0 10766 7 1 2 5158 9891
0 10767 7 1 2 5160 9892
0 10768 7 1 2 5161 8252
0 10769 5 1 1 5164
0 10770 6 1 2 5194 9245
0 10771 5 1 1 5195
0 10772 6 1 2 5214 9246
0 10773 5 1 1 5215
0 10774 6 1 2 5216 9247
0 10775 5 1 1 5217
0 10776 6 1 2 5218 9248
0 10778 3 2 2 10730 10587
0 10781 3 2 2 10731 10588
0 10784 5 4 1 5163
0 10789 6 2 2 10737 10672
0 10792 6 2 2 10738 10674
0 10796 5 1 1 5219
0 10797 6 1 2 5220 8633
0 10798 5 1 1 5221
0 10799 6 1 2 5222 8638
0 10800 6 2 2 10746 10682
0 10803 6 2 2 10747 10684
0 10806 6 2 2 10748 10686
0 10809 6 2 2 10749 10688
0 10812 6 2 2 10750 10690
0 10815 5 1 1 5223
0 10816 6 1 2 5224 9866
0 10817 6 2 2 10753 10695
0 10820 6 2 2 10754 10697
0 10823 5 1 1 5225
0 10824 6 1 2 5226 9505
0 10825 5 1 1 5227
0 10826 6 1 2 5228 9514
3 10827 6 0 2 10764 10720
0 10832 6 1 2 4281 10769
0 10833 6 1 2 4283 10771
0 10834 6 1 2 4285 10773
0 10835 6 1 2 4287 10775
0 10836 5 1 1 5229
3 10837 1 0 1 5231
3 10838 1 0 1 5232
3 10839 1 0 1 5233
3 10840 1 0 1 5234
0 10845 6 1 2 4049 10796
0 10846 6 1 2 4057 10798
0 10857 6 1 2 4686 10815
0 10862 6 1 2 4382 10823
0 10863 6 1 2 4394 10825
0 10864 7 1 2 10023 5235
0 10865 7 1 2 10024 5236
0 10866 7 1 2 9739 5237
0 10867 7 1 2 3722 5238
3 10868 6 0 2 10832 10770
3 10869 6 0 2 10833 10772
3 10870 6 0 2 10834 10774
3 10871 6 0 2 10835 10776
0 10872 5 1 1 5239
0 10873 6 1 2 5240 8616
0 10874 5 1 1 5241
0 10875 6 1 2 5242 8625
0 10876 6 2 2 10845 10797
0 10879 6 2 2 10846 10799
0 10882 5 1 1 5243
0 10883 6 1 2 5244 8645
0 10884 5 1 1 5245
0 10885 6 1 2 5246 8654
0 10886 5 1 1 5247
0 10887 6 1 2 5248 9455
0 10888 5 1 1 5249
0 10889 6 1 2 5250 9460
0 10890 5 1 1 5251
0 10891 6 1 2 5252 9862
0 10892 6 2 2 10857 10816
0 10895 5 1 1 5253
0 10896 6 1 2 5254 9494
0 10897 5 1 1 5255
0 10898 6 1 2 5256 9499
0 10899 6 2 2 10862 10824
0 10902 6 2 2 10863 10826
3 10905 3 0 2 10864 10765
3 10906 3 0 2 10865 10766
3 10907 3 0 2 10866 10767
3 10908 3 0 2 10867 10768
0 10909 6 1 2 4029 10872
0 10910 6 1 2 4041 10874
0 10915 6 1 2 4065 10882
0 10916 6 1 2 4077 10884
0 10917 6 1 2 4316 10886
0 10918 6 1 2 4324 10888
0 10919 6 1 2 4684 10890
0 10922 6 1 2 4368 10895
0 10923 6 1 2 4376 10897
0 10928 6 2 2 10909 10873
0 10931 6 2 2 10910 10875
0 10934 5 1 1 5257
0 10935 6 1 2 5258 8634
0 10936 5 1 1 5259
0 10937 6 1 2 5260 8639
0 10938 6 2 2 10915 10883
0 10941 6 2 2 10916 10885
0 10944 6 2 2 10917 10887
0 10947 6 2 2 10918 10889
0 10950 6 2 2 10919 10891
0 10953 5 1 1 5261
0 10954 6 1 2 5262 9476
0 10955 6 2 2 10922 10896
0 10958 6 2 2 10923 10898
0 10961 5 1 1 5263
0 10962 6 1 2 5264 9506
0 10963 5 1 1 5265
0 10964 6 1 2 5266 9515
0 10969 6 1 2 4051 10934
0 10970 6 1 2 4059 10936
0 10981 6 1 2 4344 10953
0 10986 6 1 2 4384 10961
0 10987 6 1 2 4396 10963
0 10988 5 1 1 5267
0 10989 6 1 2 5268 8617
0 10990 5 1 1 5269
0 10991 6 1 2 5270 8626
0 10992 6 2 2 10969 10935
0 10995 6 2 2 10970 10937
0 10998 5 1 1 5271
0 10999 6 1 2 5272 8646
0 11000 5 1 1 5273
0 11001 6 1 2 5274 8655
0 11002 5 1 1 5275
0 11003 6 1 2 5276 9456
0 11004 5 1 1 5277
0 11005 6 1 2 5278 9461
0 11006 5 1 1 5279
0 11007 6 1 2 5280 9465
0 11008 6 2 2 10981 10954
0 11011 5 1 1 5281
0 11012 6 1 2 5282 9495
0 11013 5 1 1 5301
0 11014 6 1 2 5302 9500
0 11015 6 2 2 10986 10962
0 11018 6 2 2 10987 10964
0 11023 6 1 2 4031 10988
0 11024 6 1 2 4043 10990
0 11027 6 1 2 4067 10998
0 11028 6 1 2 4079 11000
0 11029 6 1 2 4318 11002
0 11030 6 1 2 4328 11004
0 11031 6 1 2 4332 11006
0 11034 6 1 2 4370 11011
0 11035 6 1 2 4378 11013
0 11040 5 1 1 5303
0 11041 6 1 2 5304 8294
0 11042 5 1 1 5305
0 11043 6 1 2 5306 8295
0 11044 6 2 2 11023 10989
0 11047 6 2 2 11024 10991
0 11050 6 2 2 11027 10999
0 11053 6 2 2 11028 11001
0 11056 6 2 2 11029 11003
0 11059 6 2 2 11030 11005
0 11062 6 2 2 11031 11007
0 11065 5 1 1 5307
0 11066 6 1 2 5308 9477
0 11067 6 2 2 11034 11012
0 11070 6 2 2 11035 11014
0 11073 5 1 1 5309
0 11074 6 1 2 5310 9507
0 11075 5 1 1 5311
0 11076 6 1 2 5312 9516
0 11077 6 1 2 4053 11040
0 11078 6 1 2 4061 11042
0 11095 6 1 2 4346 11065
0 11098 6 1 2 4386 11073
0 11099 6 1 2 4398 11075
0 11100 6 2 2 11077 11041
0 11103 6 2 2 11078 11043
0 11106 5 1 1 5332
0 11107 6 1 2 5333 9319
0 11108 5 1 1 5334
0 11109 6 1 2 5335 9320
0 11110 5 1 1 5338
0 11111 6 1 2 5339 9381
0 11112 5 1 1 5340
0 11113 6 1 2 5341 9382
0 11114 5 1 1 5313
0 11115 6 1 2 5325 8618
0 11116 5 1 1 5326
0 11117 6 1 2 5327 8619
0 11118 5 1 1 5328
0 11119 6 1 2 5329 8647
0 11120 5 1 1 5330
0 11121 6 1 2 5331 8648
0 11122 5 1 1 5336
0 11123 6 1 2 5337 9466
0 11124 6 2 2 11095 11066
0 11127 6 2 2 11098 11074
0 11130 6 2 2 11099 11076
0 11137 6 1 2 4320 11106
0 11138 6 1 2 4330 11108
0 11139 6 1 2 4372 11110
0 11140 6 1 2 4380 11112
0 11141 6 1 2 4033 11114
0 11142 6 1 2 4045 11116
0 11143 6 1 2 4069 11118
0 11144 6 1 2 4081 11120
0 11145 6 1 2 4336 11122
0 11152 7 1 3 5344 4407 4993
0 11153 7 1 3 5342 4127 4995
0 11154 7 1 3 5345 4713 4930
0 11155 7 1 3 5343 9917 4932
0 11156 6 2 2 11137 11107
0 11159 6 2 2 11138 11109
0 11162 6 2 2 11139 11111
0 11165 6 2 2 11140 11113
0 11168 6 2 2 11141 11115
0 11171 6 2 2 11142 11117
0 11174 6 2 2 11143 11119
0 11177 6 2 2 11144 11121
0 11180 6 2 2 11145 11123
0 11183 5 1 1 5346
0 11184 6 1 2 5347 9468
0 11185 5 1 1 5348
0 11186 6 1 2 5349 9508
0 11187 5 1 1 5350
0 11188 6 1 2 5351 9509
0 11205 3 2 4 11152 11153 11154 11155
0 11210 6 1 2 4348 11183
0 11211 6 1 2 4388 11185
0 11212 6 1 2 4400 11187
0 11213 5 1 1 5360
0 11214 6 1 2 5361 8260
0 11215 5 1 1 5362
0 11216 6 1 2 5368 8261
0 11217 5 1 1 5369
0 11218 6 1 2 5370 8296
0 11219 5 1 1 5371
0 11220 6 1 2 5372 8297
0 11222 7 1 3 5354 4716 792
0 11223 7 1 3 5352 4422 793
0 11224 7 1 3 5355 4882 542
0 11225 7 1 3 5353 10132 544
0 11226 7 1 3 5358 4720 5108
0 11227 7 1 3 5356 4439 5109
0 11228 7 1 3 5359 4885 5002
0 11229 7 1 3 5357 10160 5004
0 11231 5 1 1 5373
0 11232 6 1 2 5374 9467
0 11233 6 2 2 11210 11184
0 11236 6 2 2 11211 11186
0 11239 6 2 2 11212 11188
0 11242 6 1 2 4035 11213
0 11243 6 1 2 4037 11215
0 11244 6 1 2 4071 11217
0 11245 6 1 2 4073 11219
0 11246 5 1 1 5375
0 11250 6 1 2 4338 11231
0 11252 3 2 4 11222 11223 11224 11225
0 11257 3 2 4 11226 11227 11228 11229
0 11260 6 1 2 11242 11214
0 11261 6 1 2 11243 11216
0 11262 6 1 2 11244 11218
0 11263 6 1 2 11245 11220
0 11264 5 1 1 5377
0 11265 6 1 2 5378 9322
0 11267 5 1 1 5379
0 11268 6 1 2 5380 9383
0 11269 5 1 1 5381
0 11270 6 1 2 5382 9384
0 11272 6 2 2 11250 11232
0 11277 5 1 1 11261
0 11278 7 1 2 4992 11260
0 11279 5 1 1 11263
0 11280 7 1 2 4933 11262
0 11282 6 1 2 4342 11264
0 11283 5 1 1 5383
0 11284 6 1 2 4390 11267
0 11285 6 1 2 4392 11269
0 11286 5 1 1 5385
0 11288 7 1 2 11277 5106
0 11289 7 1 2 11279 4996
0 11290 5 1 1 5387
0 11291 6 1 2 5388 9321
0 11292 6 1 2 11282 11265
0 11293 6 1 2 11284 11268
0 11294 6 1 2 11285 11270
0 11295 6 1 2 4340 11290
0 11296 5 1 1 11292
0 11297 5 1 1 11294
0 11298 7 1 2 5005 11293
0 11299 3 2 2 11288 11278
0 11302 3 2 2 11289 11280
0 11307 6 1 2 11295 11291
0 11308 7 1 2 11296 795
0 11309 7 1 2 11297 5115
0 11312 6 1 2 5391 11246
0 11313 6 1 2 5389 10836
0 11314 5 1 1 5390
0 11315 5 1 1 5392
0 11316 7 1 2 546 11307
0 11317 3 2 2 11309 11298
0 11320 6 1 2 5376 11315
0 11321 6 1 2 5230 11314
0 11323 3 2 2 11308 11316
0 11327 6 1 2 11312 11320
0 11328 6 1 2 11313 11321
0 11329 6 1 2 5393 11286
0 11331 5 1 1 5394
3 11333 5 0 1 11327
3 11334 5 0 1 11328
0 11335 6 1 2 5386 11331
0 11336 6 1 2 5395 11283
0 11337 5 1 1 5396
0 11338 6 1 2 11329 11335
0 11339 6 1 2 5384 11337
3 11340 5 0 1 11338
0 11341 6 1 2 11336 11339
3 11342 5 0 1 11341
2 2 1 1
2 3 1 1
2 4 1 1
2 6 1 5
2 7 1 5
2 8 1 5
2 10 1 9
2 11 1 9
2 13 1 12
2 14 1 12
2 16 1 15
2 17 1 15
2 19 1 18
2 20 1 18
2 21 1 18
2 22 1 18
2 24 1 23
2 25 1 23
2 27 1 26
2 28 1 26
2 30 1 29
2 31 1 29
2 33 1 32
2 34 1 32
2 36 1 35
2 37 1 35
2 39 1 38
2 40 1 38
2 42 1 41
2 43 1 41
2 45 1 44
2 46 1 44
2 48 1 47
2 49 1 47
2 51 1 50
2 52 1 50
2 67 1 66
2 68 1 66
2 71 1 70
2 72 1 70
2 90 1 89
2 91 1 89
2 92 1 89
2 93 1 89
2 95 1 94
2 96 1 94
2 98 1 97
2 99 1 97
2 101 1 100
2 102 1 100
2 104 1 103
2 105 1 103
2 107 1 106
2 108 1 106
2 116 1 115
2 117 1 115
2 119 1 118
2 120 1 118
2 122 1 121
2 123 1 121
2 125 1 124
2 126 1 124
2 128 1 127
2 129 1 127
2 131 1 130
2 132 1 130
2 136 1 135
2 137 1 135
2 139 1 138
2 140 1 138
2 142 1 141
2 143 1 141
2 145 1 144
2 146 1 144
2 148 1 147
2 149 1 147
2 243 1 242
2 244 1 242
2 246 1 245
2 247 1 245
2 249 1 248
2 250 1 248
2 252 1 251
2 253 1 251
2 255 1 254
2 256 1 254
2 258 1 257
2 259 1 257
2 261 1 260
2 262 1 260
2 264 1 263
2 265 1 263
2 266 1 263
2 268 1 267
2 269 1 267
2 270 1 267
2 272 1 271
2 273 1 271
2 275 1 274
2 276 1 274
2 278 1 277
2 279 1 277
2 281 1 280
2 282 1 280
2 284 1 283
2 285 1 283
2 287 1 286
2 288 1 286
2 290 1 289
2 291 1 289
2 292 1 289
2 294 1 293
2 295 1 293
2 297 1 296
2 298 1 296
2 300 1 299
2 301 1 299
2 302 1 299
2 304 1 303
2 305 1 303
2 306 1 303
2 308 1 307
2 309 1 307
2 311 1 310
2 312 1 310
2 314 1 313
2 315 1 313
2 317 1 316
2 318 1 316
2 320 1 319
2 321 1 319
2 323 1 322
2 324 1 322
2 326 1 325
2 327 1 325
2 329 1 328
2 330 1 328
2 332 1 331
2 333 1 331
2 335 1 334
2 336 1 334
2 338 1 337
2 339 1 337
2 341 1 340
2 342 1 340
2 344 1 343
2 345 1 343
2 347 1 346
2 348 1 346
2 350 1 349
2 351 1 349
2 353 1 352
2 354 1 352
2 356 1 355
2 357 1 355
2 359 1 358
2 360 1 358
2 362 1 361
2 363 1 361
2 365 1 364
2 366 1 364
2 368 1 367
2 369 1 367
2 370 1 367
2 371 1 367
2 372 1 367
2 373 1 367
2 374 1 367
2 375 1 367
2 376 1 367
2 377 1 367
2 378 1 367
2 379 1 367
2 380 1 367
2 381 1 367
2 383 1 382
2 384 1 382
2 385 1 382
2 386 1 382
2 389 1 469
2 390 1 469
2 391 1 494
2 392 1 494
2 393 1 528
2 394 1 528
2 395 1 575
2 396 1 575
2 397 1 578
2 398 1 578
2 399 1 590
2 400 1 590
2 401 1 593
2 402 1 593
2 403 1 596
2 404 1 596
2 405 1 599
2 406 1 599
2 407 1 599
2 408 1 599
2 409 1 604
2 410 1 604
2 411 1 604
2 412 1 604
2 413 1 609
2 414 1 609
2 415 1 609
2 416 1 609
2 417 1 614
2 418 1 614
2 419 1 614
2 420 1 614
2 421 1 614
2 422 1 614
2 423 1 614
2 424 1 614
2 425 1 614
2 426 1 614
2 427 1 625
2 428 1 625
2 429 1 628
2 430 1 628
2 431 1 628
2 432 1 632
2 433 1 632
2 434 1 632
2 435 1 636
2 436 1 636
2 437 1 636
2 438 1 636
2 439 1 644
2 440 1 644
2 441 1 644
2 442 1 644
2 443 1 644
2 444 1 644
2 445 1 651
2 446 1 651
2 447 1 651
2 448 1 651
2 449 1 651
2 450 1 657
2 451 1 657
2 452 1 660
2 453 1 660
2 454 1 660
2 455 1 660
2 456 1 660
2 457 1 666
2 458 1 666
2 459 1 666
2 460 1 666
2 461 1 666
2 462 1 676
2 463 1 676
2 464 1 676
2 465 1 676
2 466 1 676
2 468 1 682
2 470 1 682
2 471 1 682
2 472 1 682
2 473 1 682
2 474 1 689
2 475 1 689
2 476 1 689
2 477 1 689
2 479 1 689
2 480 1 695
2 481 1 695
2 483 1 695
2 485 1 695
2 487 1 700
2 488 1 700
2 490 1 700
2 491 1 700
2 493 1 708
2 495 1 708
2 496 1 708
2 497 1 708
2 498 1 708
2 499 1 708
2 500 1 715
2 502 1 715
2 503 1 715
2 504 1 715
2 506 1 715
2 508 1 721
2 510 1 721
2 512 1 721
2 514 1 721
2 516 1 721
2 518 1 727
2 520 1 727
2 521 1 727
2 522 1 727
2 523 1 727
2 524 1 734
2 525 1 734
2 526 1 734
2 527 1 734
2 529 1 734
2 530 1 734
2 531 1 734
2 532 1 742
2 533 1 742
2 534 1 742
2 536 1 742
2 538 1 742
2 540 1 750
2 542 1 750
2 544 1 750
2 546 1 750
2 548 1 759
2 550 1 759
2 552 1 762
2 554 1 762
2 555 1 762
2 557 1 762
2 558 1 762
2 560 1 768
2 562 1 768
2 564 1 768
2 566 1 768
2 568 1 768
2 570 1 774
2 572 1 774
2 574 1 774
2 576 1 774
2 577 1 774
2 579 1 780
2 580 1 780
2 581 1 780
2 583 1 780
2 584 1 780
2 586 1 786
2 587 1 786
2 588 1 786
2 589 1 786
2 591 1 786
2 592 1 786
2 594 1 786
2 595 1 794
2 597 1 794
2 598 1 794
2 600 1 794
2 601 1 794
2 602 1 800
2 603 1 800
2 605 1 800
2 606 1 800
2 607 1 800
2 608 1 806
2 610 1 806
2 611 1 806
2 612 1 806
2 613 1 806
2 615 1 814
2 616 1 814
2 617 1 814
2 618 1 814
2 619 1 814
2 620 1 814
2 621 1 821
2 622 1 821
2 623 1 821
2 624 1 821
2 626 1 821
2 627 1 827
2 629 1 827
2 630 1 827
2 631 1 827
2 633 1 827
2 634 1 833
2 635 1 833
2 637 1 833
2 638 1 833
2 639 1 833
2 640 1 839
2 645 1 839
2 646 1 839
2 647 1 839
2 648 1 839
2 649 1 845
2 650 1 845
2 652 1 845
2 653 1 845
2 654 1 845
2 655 1 845
2 656 1 845
2 658 1 853
2 659 1 853
2 661 1 853
2 662 1 853
2 663 1 853
2 664 1 859
2 665 1 859
2 667 1 859
2 668 1 859
2 669 1 859
2 670 1 865
2 671 1 865
2 675 1 865
2 677 1 865
2 678 1 865
2 679 1 871
2 680 1 871
2 681 1 957
2 683 1 957
2 684 1 957
2 685 1 957
2 686 1 957
2 687 1 957
2 690 1 1029
2 691 1 1029
2 692 1 1116
2 693 1 1116
2 694 1 1119
2 696 1 1119
2 697 1 1119
2 698 1 1119
2 699 1 1119
2 701 1 1125
2 702 1 1125
2 703 1 1125
2 704 1 1125
2 709 1 1125
2 710 1 1125
2 711 1 1132
2 712 1 1132
2 713 1 1132
2 714 1 1136
2 716 1 1136
2 717 1 1136
2 718 1 1136
2 719 1 1141
2 720 1 1141
2 722 1 1141
2 723 1 1141
2 724 1 1141
2 725 1 1147
2 726 1 1147
2 728 1 1147
2 729 1 1147
2 730 1 1147
2 731 1 1147
2 732 1 1154
2 735 1 1154
2 736 1 1154
2 737 1 1154
2 738 1 1154
2 739 1 1160
2 740 1 1160
2 741 1 1160
2 743 1 1160
2 744 1 1160
2 745 1 1160
2 746 1 1167
2 747 1 1167
2 751 1 1167
2 752 1 1167
2 753 1 1175
2 754 1 1175
2 755 1 1175
2 756 1 1175
2 757 1 1175
2 760 1 1175
2 761 1 1182
2 763 1 1182
2 764 1 1182
2 765 1 1182
2 766 1 1182
2 767 1 1182
2 769 1 1189
2 770 1 1189
2 771 1 1189
2 772 1 1189
2 773 1 1194
2 775 1 1194
2 776 1 1194
2 777 1 1194
2 778 1 1199
2 779 1 1199
2 781 1 1206
2 782 1 1206
2 783 1 1206
2 784 1 1206
2 785 1 1211
2 787 1 1211
2 788 1 1211
2 789 1 1211
2 790 1 1211
2 791 1 1211
2 792 1 1218
2 793 1 1218
2 795 1 1218
2 796 1 1222
2 797 1 1222
2 798 1 1227
2 799 1 1227
2 801 1 1227
2 802 1 1227
2 803 1 1227
2 804 1 1233
2 805 1 1233
2 807 1 1233
2 808 1 1233
2 809 1 1233
2 810 1 1233
2 811 1 1240
2 815 1 1240
2 816 1 1240
2 817 1 1244
2 818 1 1244
2 819 1 1244
2 820 1 1244
2 822 1 1249
2 823 1 1249
2 824 1 1249
2 825 1 1249
2 826 1 1249
2 828 1 1249
2 829 1 1256
2 830 1 1256
2 831 1 1256
2 832 1 1256
2 834 1 1256
2 835 1 1256
2 836 1 1263
2 837 1 1263
2 838 1 1263
2 840 1 1263
2 841 1 1263
2 842 1 1263
2 843 1 1270
2 844 1 1270
2 846 1 1270
2 847 1 1270
2 848 1 1270
2 849 1 1270
2 850 1 1277
2 851 1 1277
2 852 1 1277
2 854 1 1277
2 855 1 1277
2 856 1 1277
2 857 1 1284
2 858 1 1284
2 860 1 1287
2 861 1 1287
2 862 1 1290
2 863 1 1290
2 864 1 1293
2 866 1 1293
2 867 1 1296
2 868 1 1296
2 869 1 1299
2 870 1 1299
2 872 1 1302
2 873 1 1302
2 874 1 1305
2 875 1 1305
2 876 1 1308
2 877 1 1308
2 878 1 1311
2 879 1 1311
2 880 1 1314
2 888 1 1314
2 890 1 1317
2 891 1 1317
2 892 1 1320
2 893 1 1320
2 894 1 1323
2 895 1 1323
2 896 1 1326
2 897 1 1326
2 898 1 1329
2 899 1 1329
2 900 1 1332
2 901 1 1332
2 902 1 1335
2 903 1 1335
2 904 1 1338
2 905 1 1338
2 906 1 1341
2 907 1 1341
2 908 1 1344
2 909 1 1344
2 910 1 1347
2 911 1 1347
2 912 1 1350
2 913 1 1350
2 914 1 1353
2 915 1 1353
2 916 1 1356
2 917 1 1356
2 918 1 1359
2 919 1 1359
2 920 1 1362
2 921 1 1362
2 922 1 1365
2 923 1 1365
2 924 1 1368
2 925 1 1368
2 926 1 1371
2 927 1 1371
2 928 1 1374
2 929 1 1374
2 930 1 1377
2 931 1 1377
2 932 1 1380
2 933 1 1380
2 934 1 1383
2 935 1 1383
2 936 1 1386
2 937 1 1386
2 938 1 1389
2 939 1 1389
2 940 1 1392
2 941 1 1392
2 942 1 1395
2 943 1 1395
2 944 1 1398
2 946 1 1398
2 947 1 1401
2 948 1 1401
2 949 1 1404
2 950 1 1404
2 951 1 1407
2 952 1 1407
2 953 1 1410
2 954 1 1410
2 955 1 1413
2 956 1 1413
2 958 1 1416
2 959 1 1416
2 960 1 1419
2 961 1 1419
2 962 1 1422
2 963 1 1422
2 964 1 1425
2 965 1 1425
2 966 1 1428
2 967 1 1428
2 968 1 1431
2 969 1 1431
2 970 1 1434
2 971 1 1434
2 972 1 1437
2 973 1 1437
2 974 1 1440
2 975 1 1440
2 976 1 1443
2 977 1 1443
2 978 1 1446
2 979 1 1446
2 980 1 1449
2 981 1 1449
2 982 1 1452
2 983 1 1452
2 984 1 1455
2 985 1 1455
2 986 1 1458
2 987 1 1458
2 988 1 1461
2 989 1 1461
2 990 1 1464
2 991 1 1464
2 992 1 1467
2 993 1 1467
2 994 1 1470
2 995 1 1470
2 996 1 1473
2 997 1 1473
2 998 1 1476
2 999 1 1476
2 1000 1 1479
2 1001 1 1479
2 1002 1 1482
2 1003 1 1482
2 1004 1 1485
2 1005 1 1485
2 1006 1 1537
2 1007 1 1537
2 1008 1 1537
2 1009 1 1537
2 1010 1 1537
2 1011 1 1551
2 1012 1 1551
2 1013 1 1703
2 1014 1 1703
2 1015 1 1708
2 1016 1 1708
2 1017 1 1713
2 1018 1 1713
2 1019 1 1721
2 1020 1 1721
2 1021 1 1758
2 1022 1 1758
2 1023 1 1783
2 1024 1 1783
2 1025 1 1783
2 1026 1 1783
2 1027 1 1783
2 1030 1 1789
2 1031 1 1789
2 1032 1 1789
2 1033 1 1799
2 1034 1 1799
2 1035 1 1799
2 1036 1 1799
2 1037 1 1799
2 1038 1 1805
2 1039 1 1805
2 1040 1 1805
2 1041 1 1805
2 1042 1 1805
2 1043 1 1845
2 1044 1 1845
2 1045 1 1845
2 1046 1 1845
2 1047 1 1845
2 1048 1 1851
2 1049 1 1851
2 1050 1 1851
2 1051 1 1851
2 1052 1 1851
2 1053 1 1885
2 1054 1 1885
2 1055 1 1885
2 1056 1 1885
2 1057 1 1885
2 1058 1 1885
2 1059 1 1892
2 1060 1 1892
2 1061 1 1892
2 1062 1 1892
2 1063 1 1892
2 1064 1 1892
2 1065 1 1899
2 1066 1 1899
2 1067 1 1899
2 1068 1 1899
2 1069 1 1899
2 1070 1 1899
2 1071 1 1906
2 1072 1 1906
2 1073 1 1906
2 1074 1 1906
2 1075 1 1906
2 1076 1 1906
2 1077 1 1913
2 1078 1 1913
2 1079 1 1913
2 1080 1 1913
2 1081 1 1913
2 1082 1 1919
2 1083 1 1919
2 1084 1 1919
2 1085 1 1919
2 1086 1 1919
2 1087 1 1919
2 1088 1 1947
2 1089 1 1947
2 1090 1 1947
2 1091 1 1947
2 1092 1 1947
2 1093 1 1953
2 1094 1 1953
2 1095 1 1953
2 1096 1 1977
2 1097 1 1977
2 1098 1 1977
2 1099 1 1977
2 1100 1 1977
2 1101 1 1983
2 1102 1 1983
2 1103 1 1983
2 1104 1 1983
2 1105 1 1983
2 1106 1 1997
2 1107 1 1997
2 1108 1 1997
2 1117 1 1997
2 1118 1 1997
2 1120 1 2003
2 1121 1 2003
2 1122 1 2003
2 1123 1 2003
2 1124 1 2003
2 1126 1 2003
2 1127 1 2024
2 1128 1 2024
2 1129 1 2024
2 1130 1 2024
2 1131 1 2024
2 1133 1 2024
2 1134 1 2031
2 1135 1 2031
2 1137 1 2031
2 1138 1 2031
2 1139 1 2031
2 1140 1 2031
2 1142 1 2038
2 1143 1 2038
2 1144 1 2038
2 1145 1 2038
2 1146 1 2038
2 1148 1 2038
2 1149 1 2045
2 1150 1 2045
2 1151 1 2045
2 1152 1 2045
2 1153 1 2045
2 1155 1 2045
2 1156 1 2052
2 1157 1 2052
2 1158 1 2052
2 1159 1 2052
2 1161 1 2052
2 1162 1 2058
2 1163 1 2058
2 1164 1 2058
2 1165 1 2058
2 1166 1 2058
2 1168 1 2074
2 1169 1 2074
2 1170 1 2081
2 1171 1 2081
2 1172 1 2086
2 1173 1 2086
2 1176 1 2231
2 1177 1 2231
2 1178 1 2235
2 1179 1 2235
2 1180 1 2257
2 1181 1 2257
2 1183 1 2257
2 1184 1 2257
2 1185 1 2257
2 1186 1 2257
2 1187 1 2257
2 1188 1 2257
2 1190 1 2257
2 1191 1 2269
2 1192 1 2269
2 1193 1 2269
2 1195 1 2269
2 1196 1 2287
2 1197 1 2287
2 1198 1 2287
2 1200 1 2287
2 1201 1 2287
2 1202 1 2293
2 1203 1 2293
2 1204 1 2293
2 1205 1 2293
2 1207 1 2293
2 1208 1 2309
2 1209 1 2309
2 1210 1 2309
2 1212 1 2309
2 1213 1 2309
2 1214 1 2315
2 1215 1 2315
2 1216 1 2315
2 1217 1 2315
2 1219 1 2315
2 1220 1 2331
2 1221 1 2331
2 1223 1 2331
2 1224 1 2331
2 1225 1 2331
2 1226 1 2368
2 1228 1 2368
2 1229 1 2368
2 1230 1 2368
2 1231 1 2368
2 1232 1 2384
2 1234 1 2384
2 1235 1 2384
2 1236 1 2384
2 1237 1 2384
2 1238 1 2390
2 1239 1 2390
2 1241 1 2390
2 1242 1 2390
2 1243 1 2390
2 1245 1 2406
2 1246 1 2406
2 1247 1 2406
2 1248 1 2406
2 1250 1 2406
2 1251 1 2412
2 1252 1 2412
2 1253 1 2412
2 1254 1 2412
2 1255 1 2412
2 1257 1 2442
2 1258 1 2442
2 1259 1 2442
2 1260 1 2446
2 1261 1 2446
2 1262 1 2446
2 1264 1 2450
2 1265 1 2450
2 1266 1 2450
2 1267 1 2454
2 1268 1 2454
2 1269 1 2454
2 1271 1 2458
2 1272 1 2458
2 1273 1 2458
2 1274 1 2462
2 1275 1 2462
2 1276 1 2462
2 1278 1 2466
2 1279 1 2466
2 1280 1 2466
2 1281 1 2470
2 1282 1 2470
2 1283 1 2470
2 1285 1 2474
2 1286 1 2474
2 1288 1 2474
2 1289 1 2478
2 1291 1 2478
2 1292 1 2478
2 1294 1 2482
2 1295 1 2482
2 1297 1 2482
2 1298 1 2482
2 1300 1 2482
2 1301 1 2488
2 1303 1 2488
2 1304 1 2488
2 1306 1 2488
2 1307 1 2488
2 1309 1 2488
2 1310 1 2488
2 1312 1 2496
2 1313 1 2496
2 1315 1 2496
2 1316 1 2496
2 1318 1 2496
2 1319 1 2502
2 1321 1 2502
2 1322 1 2502
2 1324 1 2502
2 1325 1 2502
2 1327 1 2508
2 1328 1 2508
2 1330 1 2508
2 1331 1 2508
2 1333 1 2508
2 1334 1 2523
2 1336 1 2523
2 1337 1 2523
2 1339 1 2523
2 1340 1 2523
2 1342 1 2533
2 1343 1 2533
2 1345 1 2533
2 1346 1 2538
2 1348 1 2538
2 1349 1 2538
2 1351 1 2542
2 1352 1 2542
2 1354 1 2542
2 1355 1 2546
2 1357 1 2546
2 1358 1 2546
2 1360 1 2550
2 1361 1 2550
2 1363 1 2550
2 1364 1 2554
2 1366 1 2554
2 1367 1 2554
2 1369 1 2554
2 1370 1 2554
2 1372 1 2554
2 1373 1 2561
2 1375 1 2561
2 1376 1 2561
2 1378 1 2561
2 1379 1 2561
2 1381 1 2567
2 1382 1 2567
2 1384 1 2567
2 1385 1 2567
2 1387 1 2567
2 1388 1 2573
2 1390 1 2573
2 1391 1 2573
2 1393 1 2573
2 1394 1 2573
2 1396 1 2604
2 1397 1 2604
2 1399 1 2607
2 1400 1 2607
2 1402 1 2607
2 1403 1 2611
2 1405 1 2611
2 1406 1 2611
2 1408 1 2615
2 1409 1 2615
2 1411 1 2615
2 1412 1 2619
2 1414 1 2619
2 1415 1 2619
2 1417 1 2619
2 1418 1 2619
2 1420 1 2619
2 1421 1 2626
2 1423 1 2626
2 1424 1 2626
2 1426 1 2626
2 1427 1 2626
2 1429 1 2632
2 1430 1 2632
2 1432 1 2632
2 1433 1 2632
2 1435 1 2632
2 1436 1 2638
2 1438 1 2638
2 1439 1 2638
2 1441 1 2638
2 1442 1 2638
2 1444 1 2644
2 1445 1 2644
2 1447 1 2644
2 1448 1 2644
2 1450 1 2644
2 1451 1 2650
2 1453 1 2650
2 1454 1 2654
2 1456 1 2654
2 1457 1 2654
2 1459 1 2658
2 1460 1 2658
2 1462 1 2658
2 1463 1 2662
2 1465 1 2662
2 1466 1 2662
2 1468 1 2666
2 1469 1 2666
2 1471 1 2666
2 1472 1 2670
2 1474 1 2670
2 1475 1 2670
2 1477 1 2674
2 1478 1 2674
2 1480 1 2674
2 1481 1 2674
2 1483 1 2674
2 1484 1 2680
2 1486 1 2680
2 1487 1 2688
2 1488 1 2688
2 1491 1 2688
2 1492 1 2692
2 1493 1 2692
2 1494 1 2692
2 1495 1 2696
2 1496 1 2696
2 1497 1 2696
2 1498 1 2700
2 1499 1 2700
2 1500 1 2700
2 1501 1 2704
2 1502 1 2704
2 1503 1 2704
2 1504 1 2729
2 1505 1 2729
2 1506 1 2729
2 1507 1 2733
2 1508 1 2733
2 1509 1 2733
2 1510 1 2737
2 1511 1 2737
2 1512 1 2737
2 1513 1 2741
2 1514 1 2741
2 1515 1 2741
2 1516 1 2745
2 1517 1 2745
2 1518 1 2745
2 1519 1 2749
2 1520 1 2749
2 1521 1 2749
2 1522 1 2753
2 1523 1 2753
2 1524 1 2753
2 1525 1 2757
2 1526 1 2757
2 1527 1 2757
2 1528 1 2761
2 1529 1 2761
2 1530 1 2761
2 1531 1 2766
2 1532 1 2766
2 1533 1 2769
2 1534 1 2769
2 1535 1 2772
2 1536 1 2772
2 1538 1 2775
2 1539 1 2775
2 1540 1 2778
2 1541 1 2778
2 1542 1 2781
2 1543 1 2781
2 1544 1 2784
2 1545 1 2784
2 1546 1 2787
2 1547 1 2787
2 1548 1 2790
2 1549 1 2790
2 1550 1 2793
2 1552 1 2793
2 1553 1 2796
2 1554 1 2796
2 1555 1 3061
2 1556 1 3061
2 1557 1 3064
2 1558 1 3064
2 1559 1 3067
2 1560 1 3067
2 1561 1 3070
2 1562 1 3070
2 1563 1 3073
2 1564 1 3073
2 1565 1 3080
2 1566 1 3080
2 1567 1 3097
2 1568 1 3097
2 1569 1 3097
2 1570 1 3101
2 1571 1 3101
2 1572 1 3101
2 1573 1 3101
2 1574 1 3101
2 1575 1 3107
2 1576 1 3107
2 1577 1 3107
2 1578 1 3107
2 1579 1 3107
2 1580 1 3107
2 1581 1 3114
2 1582 1 3114
2 1583 1 3114
2 1584 1 3114
2 1585 1 3114
2 1586 1 3114
2 1587 1 3114
2 1588 1 3122
2 1589 1 3122
2 1590 1 3122
2 1591 1 3126
2 1592 1 3126
2 1593 1 3126
2 1594 1 3131
2 1595 1 3131
2 1596 1 3137
2 1597 1 3137
2 1598 1 3140
2 1599 1 3140
2 1600 1 3140
2 1601 1 3144
2 1602 1 3144
2 1603 1 3144
2 1604 1 3144
2 1605 1 3149
2 1606 1 3149
2 1607 1 3149
2 1608 1 3149
2 1609 1 3149
2 1610 1 3155
2 1611 1 3155
2 1612 1 3155
2 1613 1 3159
2 1614 1 3159
2 1615 1 3159
2 1616 1 3169
2 1617 1 3169
2 1618 1 3169
2 1619 1 3173
2 1620 1 3173
2 1621 1 3173
2 1622 1 3173
2 1623 1 3178
2 1624 1 3178
2 1625 1 3178
2 1626 1 3178
2 1627 1 3178
2 1628 1 3185
2 1629 1 3185
2 1630 1 3185
2 1631 1 3189
2 1632 1 3189
2 1633 1 3189
2 1634 1 3189
2 1635 1 3189
2 1636 1 3195
2 1637 1 3195
2 1638 1 3195
2 1639 1 3195
2 1640 1 3195
2 1641 1 3195
2 1642 1 3202
2 1643 1 3202
2 1644 1 3202
2 1645 1 3202
2 1646 1 3202
2 1647 1 3202
2 1648 1 3202
2 1650 1 3211
2 1651 1 3211
2 1652 1 3211
2 1653 1 3215
2 1654 1 3215
2 1655 1 3215
2 1656 1 3215
2 1657 1 3215
2 1658 1 3221
2 1659 1 3221
2 1660 1 3221
2 1661 1 3221
2 1662 1 3221
2 1663 1 3221
2 1664 1 3229
2 1665 1 3229
2 1666 1 3232
2 1667 1 3232
2 1668 1 3232
2 1669 1 3236
2 1670 1 3236
2 1671 1 3236
2 1672 1 3236
2 1673 1 3241
2 1674 1 3241
2 1675 1 3241
2 1676 1 3241
2 1677 1 3241
2 1678 1 3247
2 1679 1 3247
2 1680 1 3247
2 1681 1 3251
2 1682 1 3251
2 1683 1 3251
2 1684 1 3255
2 1685 1 3255
2 1686 1 3255
2 1687 1 3259
2 1688 1 3259
2 1689 1 3259
2 1690 1 3263
2 1691 1 3263
2 1692 1 3263
2 1693 1 3267
2 1694 1 3267
2 1695 1 3267
2 1696 1 3267
2 1697 1 3267
2 1698 1 3273
2 1699 1 3273
2 1700 1 3273
2 1701 1 3273
2 1702 1 3273
2 1704 1 3273
2 1705 1 3273
2 1706 1 3281
2 1707 1 3281
2 1709 1 3281
2 1710 1 3281
2 1711 1 3281
2 1712 1 3287
2 1714 1 3287
2 1715 1 3287
2 1716 1 3287
2 1717 1 3287
2 1718 1 3293
2 1719 1 3293
2 1720 1 3293
2 1722 1 3293
2 1723 1 3293
2 1724 1 3299
2 1725 1 3299
2 1726 1 3299
2 1727 1 3303
2 1728 1 3303
2 1729 1 3303
2 1730 1 3307
2 1731 1 3307
2 1732 1 3307
2 1733 1 3311
2 1734 1 3311
2 1735 1 3311
2 1736 1 3315
2 1737 1 3315
2 1738 1 3315
2 1739 1 3315
2 1740 1 3315
2 1741 1 3315
2 1742 1 3322
2 1743 1 3322
2 1744 1 3322
2 1745 1 3322
2 1746 1 3322
2 1747 1 3328
2 1748 1 3328
2 1749 1 3328
2 1750 1 3328
2 1751 1 3328
2 1752 1 3334
2 1753 1 3334
2 1754 1 3334
2 1755 1 3334
2 1756 1 3334
2 1757 1 3340
2 1759 1 3340
2 1760 1 3343
2 1761 1 3343
2 1762 1 3343
2 1763 1 3343
2 1764 1 3343
2 1765 1 3349
2 1766 1 3349
2 1767 1 3349
2 1768 1 3349
2 1769 1 3349
2 1770 1 3355
2 1771 1 3355
2 1772 1 3355
2 1773 1 3355
2 1774 1 3355
2 1775 1 3375
2 1776 1 3375
2 1777 1 3375
2 1778 1 3381
2 1779 1 3381
2 1780 1 3384
2 1784 1 3384
2 1785 1 3384
2 1786 1 3384
2 1787 1 3384
2 1788 1 3390
2 1790 1 3390
2 1791 1 3390
2 1792 1 3390
2 1800 1 3390
2 1801 1 3390
2 1802 1 3390
2 1803 1 3398
2 1804 1 3398
2 1806 1 3398
2 1807 1 3398
2 1808 1 3398
2 1809 1 3404
2 1810 1 3404
2 1823 1 3404
2 1824 1 3404
2 1825 1 3404
2 1826 1 3410
2 1827 1 3410
2 1831 1 3410
2 1836 1 3410
2 1837 1 3410
2 1838 1 3416
2 1844 1 3416
2 1846 1 3416
2 1847 1 3420
2 1848 1 3420
2 1849 1 3420
2 1850 1 3424
2 1852 1 3424
2 1853 1 3424
2 1854 1 3428
2 1855 1 3428
2 1856 1 3428
2 1886 1 3432
2 1887 1 3432
2 1888 1 3432
2 1889 1 3436
2 1890 1 3436
2 1891 1 3436
2 1893 1 3440
2 1894 1 3440
2 1895 1 3440
2 1896 1 3444
2 1897 1 3444
2 1898 1 3444
2 1900 1 3448
2 1901 1 3448
2 1902 1 3448
2 1903 1 3454
2 1904 1 3454
2 1905 1 3454
2 1907 1 3458
2 1908 1 3458
2 1909 1 3458
2 1910 1 3462
2 1911 1 3462
2 1912 1 3462
2 1914 1 3466
2 1915 1 3466
2 1916 1 3466
2 1917 1 3470
2 1918 1 3470
2 1920 1 3470
2 1921 1 3474
2 1922 1 3474
2 1923 1 3474
2 1924 1 3478
2 1925 1 3478
2 1948 1 3478
2 1949 1 3482
2 1950 1 3482
2 1951 1 3482
2 1952 1 3487
2 1954 1 3487
2 1955 1 3490
2 1956 1 3490
2 1964 1 3493
2 1978 1 3493
2 1979 1 3496
2 1980 1 3496
2 1981 1 3499
2 1982 1 3499
2 1984 1 3502
2 1985 1 3502
2 1986 1 3507
2 1987 1 3507
2 1988 1 3510
2 1998 1 3510
2 1999 1 3515
2 2000 1 3515
2 2001 1 3518
2 2002 1 3518
2 2004 1 3521
2 2005 1 3521
2 2006 1 3524
2 2007 1 3524
2 2008 1 3527
2 2009 1 3527
2 2025 1 3530
2 2026 1 3530
2 2027 1 3535
2 2028 1 3535
2 2029 1 3539
2 2030 1 3539
2 2032 1 3542
2 2033 1 3542
2 2034 1 3545
2 2035 1 3545
2 2036 1 3548
2 2037 1 3548
2 2039 1 3553
2 2040 1 3553
2 2041 1 3557
2 2042 1 3557
2 2043 1 3560
2 2044 1 3560
2 2046 1 3563
2 2047 1 3563
2 2048 1 3566
2 2049 1 3566
2 2050 1 3571
2 2051 1 3571
2 2053 1 3574
2 2054 1 3574
2 2055 1 3577
2 2056 1 3577
2 2057 1 3580
2 2059 1 3580
2 2060 1 3583
2 2061 1 3583
2 2062 1 3586
2 2063 1 3586
2 2075 1 3589
2 2076 1 3589
2 2077 1 3592
2 2078 1 3592
2 2079 1 3595
2 2080 1 3595
2 2082 1 3598
2 2083 1 3598
2 2084 1 3601
2 2085 1 3601
2 2087 1 3604
2 2088 1 3604
2 2089 1 3607
2 2090 1 3607
2 2091 1 3610
2 2092 1 3610
2 2093 1 3613
2 2094 1 3613
2 2095 1 3616
2 2096 1 3616
2 2097 1 3619
2 2098 1 3619
2 2099 1 3622
2 2100 1 3622
2 2101 1 3625
2 2102 1 3625
2 2103 1 3628
2 2104 1 3628
2 2105 1 3631
2 2106 1 3631
2 2109 1 3634
2 2116 1 3634
2 2118 1 3637
2 2119 1 3637
2 2120 1 3640
2 2121 1 3640
2 2122 1 3643
2 2123 1 3643
2 2124 1 3646
2 2125 1 3646
2 2126 1 3649
2 2127 1 3649
2 2128 1 3652
2 2129 1 3652
2 2130 1 3655
2 2131 1 3655
2 2132 1 3658
2 2133 1 3658
2 2134 1 3661
2 2135 1 3661
2 2136 1 3664
2 2137 1 3664
2 2138 1 3667
2 2139 1 3667
2 2140 1 3670
2 2141 1 3670
2 2142 1 3673
2 2143 1 3673
2 2144 1 3676
2 2145 1 3676
2 2146 1 3679
2 2147 1 3679
2 2148 1 3682
2 2149 1 3682
2 2150 1 3685
2 2151 1 3685
2 2152 1 3688
2 2153 1 3688
2 2154 1 3691
2 2155 1 3691
2 2156 1 3694
2 2157 1 3694
2 2158 1 3697
2 2159 1 3697
2 2160 1 3700
2 2161 1 3700
2 2162 1 3703
2 2163 1 3703
2 2164 1 3706
2 2165 1 3706
2 2166 1 3709
2 2167 1 3709
2 2168 1 3712
2 2169 1 3712
2 2170 1 3715
2 2173 1 3715
2 2174 1 3718
2 2175 1 3718
2 2176 1 3721
2 2177 1 3721
2 2178 1 3724
2 2179 1 3724
2 2180 1 3727
2 2181 1 3727
2 2182 1 3730
2 2183 1 3730
2 2184 1 3733
2 2185 1 3733
2 2186 1 3736
2 2187 1 3736
2 2188 1 3739
2 2189 1 3739
2 2190 1 3742
2 2191 1 3742
2 2192 1 3745
2 2193 1 3745
2 2194 1 3748
2 2195 1 3748
2 2196 1 3751
2 2197 1 3751
2 2198 1 3754
2 2199 1 3754
2 2200 1 3757
2 2201 1 3757
2 2202 1 3760
2 2203 1 3760
2 2204 1 3763
2 2205 1 3763
2 2206 1 3766
2 2207 1 3766
2 2208 1 3769
2 2209 1 3769
2 2210 1 3772
2 2211 1 3772
2 2212 1 3775
2 2213 1 3775
2 2214 1 3778
2 2215 1 3778
2 2216 1 3783
2 2217 1 3783
2 2218 1 3786
2 2219 1 3786
2 2220 1 3789
2 2221 1 3789
2 2222 1 3792
2 2223 1 3792
2 2224 1 3795
2 2225 1 3795
2 2226 1 3798
2 2227 1 3798
2 2228 1 3801
2 2229 1 3801
2 2232 1 3804
2 2233 1 3804
2 2234 1 3807
2 2236 1 3807
2 2237 1 3810
2 2238 1 3810
2 2258 1 3813
2 2259 1 3813
2 2260 1 3816
2 2261 1 3816
2 2262 1 3819
2 2263 1 3819
2 2264 1 3822
2 2265 1 3822
2 2266 1 3825
2 2270 1 3825
2 2271 1 3828
2 2272 1 3828
2 2273 1 3831
2 2276 1 3831
2 2288 1 3834
2 2289 1 3834
2 2290 1 3837
2 2291 1 3837
2 2292 1 3840
2 2294 1 3840
2 2295 1 3843
2 2296 1 3843
2 2297 1 3846
2 2298 1 3846
2 2310 1 3849
2 2311 1 3849
2 2312 1 3852
2 2313 1 3852
2 2314 1 3855
2 2316 1 3855
2 2317 1 3858
2 2318 1 3858
2 2319 1 3861
2 2320 1 3861
2 2332 1 3864
2 2333 1 3864
2 2334 1 3867
2 2335 1 3867
2 2336 1 3870
2 2369 1 3870
2 2370 1 3873
2 2371 1 3873
2 2372 1 3876
2 2373 1 3876
2 2385 1 3879
2 2386 1 3879
2 2387 1 3882
2 2388 1 3882
2 2389 1 3885
2 2391 1 3885
2 2392 1 3888
2 2393 1 3888
2 2394 1 3891
2 2395 1 3891
2 2407 1 4193
2 2408 1 4193
2 2409 1 4193
2 2410 1 4303
2 2411 1 4303
2 2413 1 4545
2 2414 1 4545
2 2415 1 4545
2 2416 1 4549
2 2417 1 4549
2 2438 1 4549
2 2439 1 4549
2 2440 1 4549
2 2443 1 4555
2 2444 1 4555
2 2445 1 4555
2 2447 1 4555
2 2448 1 4555
2 2449 1 4555
2 2451 1 4563
2 2452 1 4563
2 2453 1 4566
2 2455 1 4566
2 2456 1 4566
2 2457 1 4570
2 2459 1 4570
2 2460 1 4570
2 2461 1 4570
2 2463 1 4577
2 2464 1 4577
2 2465 1 4577
2 2467 1 4581
2 2468 1 4581
2 2469 1 4581
2 2471 1 4581
2 2472 1 4586
2 2473 1 4586
2 2475 1 4586
2 2476 1 4586
2 2477 1 4586
2 2479 1 4593
2 2480 1 4593
2 2481 1 4593
2 2483 1 4597
2 2484 1 4597
2 2485 1 4597
2 2486 1 4597
2 2487 1 4597
2 2489 1 4603
2 2490 1 4603
2 2491 1 4603
2 2492 1 4603
2 2493 1 4603
2 2494 1 4603
2 2495 1 4657
2 2497 1 4657
2 2498 1 4657
2 2499 1 4661
2 2500 1 4661
2 2501 1 4661
2 2503 1 4661
2 2504 1 4661
2 2505 1 4667
2 2506 1 4667
2 2507 1 4667
2 2509 1 4667
2 2510 1 4667
2 2511 1 4667
2 2512 1 4675
2 2513 1 4675
2 2514 1 4678
2 2515 1 4678
2 2516 1 4678
2 2517 1 4682
2 2518 1 4682
2 2519 1 4682
2 2520 1 4682
2 2521 1 4687
2 2522 1 4687
2 2524 1 4687
2 2525 1 4687
2 2526 1 4687
2 2527 1 4702
2 2528 1 4702
2 2529 1 4702
2 2530 1 4706
2 2531 1 4706
2 2532 1 4706
2 2534 1 4706
2 2535 1 4711
2 2536 1 4711
2 2539 1 4711
2 2540 1 4711
2 2541 1 4711
2 2543 1 4718
2 2544 1 4718
2 2545 1 4718
2 2547 1 4722
2 2548 1 4722
2 2549 1 4722
2 2551 1 4722
2 2552 1 4722
2 2553 1 4728
2 2555 1 4728
2 2556 1 4728
2 2557 1 4728
2 2558 1 4728
2 2559 1 4728
2 2560 1 4735
2 2562 1 4735
2 2563 1 4735
2 2564 1 4735
2 2565 1 4735
2 2566 1 4735
2 2568 1 4735
2 2569 1 4769
2 2570 1 4769
2 2571 1 4769
2 2572 1 4769
2 2574 1 4769
2 2575 1 4784
2 2576 1 4784
2 2577 1 4790
2 2578 1 4790
2 2579 1 4796
2 2580 1 4796
2 2581 1 4803
2 2582 1 4803
2 2583 1 4806
2 2584 1 4806
2 2585 1 4810
2 2586 1 4810
2 2587 1 4814
2 2588 1 4814
2 2589 1 4817
2 2590 1 4817
2 2591 1 4820
2 2592 1 4820
2 2593 1 4823
2 2594 1 4823
2 2595 1 4826
2 2596 1 4826
2 2597 1 4829
2 2598 1 4829
2 2599 1 4832
2 2600 1 4832
2 2601 1 4835
2 2602 1 4835
2 2603 1 4838
2 2605 1 4838
2 2606 1 4841
2 2608 1 4841
2 2609 1 4844
2 2610 1 4844
2 2612 1 4847
2 2613 1 4847
2 2614 1 4850
2 2616 1 4850
2 2617 1 4853
2 2618 1 4853
2 2620 1 4856
2 2621 1 4856
2 2622 1 4859
2 2623 1 4859
2 2624 1 4862
2 2625 1 4862
2 2627 1 4865
2 2628 1 4865
2 2629 1 4868
2 2630 1 4868
2 2631 1 4871
2 2633 1 4871
2 2634 1 4874
2 2635 1 4874
2 2636 1 4877
2 2637 1 4877
2 2639 1 4880
2 2640 1 4880
2 2641 1 4883
2 2642 1 4883
2 2643 1 4886
2 2645 1 4886
2 2646 1 4889
2 2647 1 4889
2 2648 1 4892
2 2649 1 4892
2 2651 1 4895
2 2652 1 4895
2 2655 1 4898
2 2656 1 4898
2 2657 1 4901
2 2659 1 4901
2 2660 1 4904
2 2661 1 4904
2 2663 1 4907
2 2664 1 4907
2 2665 1 4910
2 2667 1 4910
2 2668 1 4913
2 2669 1 4913
2 2671 1 4916
2 2672 1 4916
2 2673 1 4919
2 2675 1 4919
2 2676 1 4922
2 2677 1 4922
2 2678 1 4925
2 2679 1 4925
2 2681 1 4928
2 2682 1 4928
2 2683 1 4931
2 2684 1 4931
2 2685 1 4934
2 2686 1 4934
2 2687 1 4937
2 2689 1 4937
2 2690 1 4940
2 2691 1 4940
2 2693 1 4943
2 2694 1 4943
2 2695 1 4946
2 2697 1 4946
2 2698 1 4949
2 2699 1 4949
2 2701 1 4952
2 2702 1 4952
2 2703 1 4955
2 2705 1 4955
2 2706 1 4958
2 2707 1 4958
2 2708 1 4961
2 2709 1 4961
2 2710 1 4964
2 2711 1 4964
2 2712 1 4967
2 2713 1 4967
2 2714 1 4970
2 2715 1 4970
2 2716 1 4973
2 2717 1 4973
2 2718 1 4976
2 2719 1 4976
2 2720 1 4979
2 2721 1 4979
2 2722 1 4982
2 2723 1 4982
2 2724 1 4985
2 2725 1 4985
2 2726 1 4988
2 2727 1 4988
2 2730 1 4991
2 2731 1 4991
2 2732 1 4994
2 2734 1 4994
2 2735 1 4997
2 2736 1 4997
2 2738 1 5000
2 2739 1 5000
2 2740 1 5003
2 2742 1 5003
2 2743 1 5006
2 2744 1 5006
2 2746 1 5009
2 2747 1 5009
2 2748 1 5012
2 2750 1 5012
2 2751 1 5015
2 2752 1 5015
2 2754 1 5018
2 2755 1 5018
2 2756 1 5021
2 2758 1 5021
2 2759 1 5024
2 2760 1 5024
2 2762 1 5027
2 2763 1 5027
2 2764 1 5030
2 2767 1 5030
2 2768 1 5033
2 2770 1 5033
2 2771 1 5036
2 2773 1 5036
2 2774 1 5039
2 2776 1 5039
2 2777 1 5042
2 2779 1 5042
2 2780 1 5049
2 2782 1 5049
2 2783 1 5052
2 2785 1 5052
2 2786 1 5055
2 2788 1 5055
2 2789 1 5058
2 2791 1 5058
2 2792 1 5061
2 2794 1 5061
2 2795 1 5068
2 2797 1 5068
2 2798 1 5071
2 2799 1 5071
2 2800 1 5074
2 2801 1 5074
2 2802 1 5077
2 2803 1 5077
2 2804 1 5080
2 2805 1 5080
2 2806 1 5083
2 2807 1 5083
2 2808 1 5086
2 2809 1 5086
2 2810 1 5089
2 2811 1 5089
2 2812 1 5092
2 2813 1 5092
2 2814 1 5095
2 2815 1 5095
2 2816 1 5098
2 2817 1 5098
2 2818 1 5101
2 2819 1 5101
2 2820 1 5104
2 2821 1 5104
2 2822 1 5107
2 2823 1 5107
2 2824 1 5114
2 2825 1 5114
2 2826 1 5117
2 2827 1 5117
2 2828 1 5120
2 2829 1 5120
2 2830 1 5123
2 2831 1 5123
2 2832 1 5126
2 2833 1 5126
2 2834 1 5129
2 2835 1 5129
2 2836 1 5132
2 2837 1 5132
2 2838 1 5135
2 2839 1 5135
2 2840 1 5138
2 2841 1 5138
2 2842 1 5141
2 2843 1 5141
2 2844 1 5144
2 2845 1 5144
2 2846 1 5147
2 2847 1 5147
2 2848 1 5150
2 2849 1 5150
2 2850 1 5153
2 2851 1 5153
2 2852 1 5156
2 2853 1 5156
2 2854 1 5159
2 2855 1 5159
2 2856 1 5162
2 2857 1 5162
2 2858 1 5632
2 2859 1 5632
2 2860 1 5632
2 2861 1 5632
2 2862 1 5632
2 2863 1 5632
2 2864 1 5632
2 2865 1 5640
2 2870 1 5640
2 2871 1 5640
2 2872 1 5640
2 2873 1 5640
2 2874 1 5640
2 2875 1 5640
2 2876 1 5640
2 2877 1 5640
2 2879 1 5640
2 2880 1 5640
2 2881 1 5640
2 2882 1 5640
2 2883 1 5654
2 2884 1 5654
2 2885 1 5654
2 2886 1 5654
2 2887 1 5654
2 2888 1 5654
2 2889 1 5654
2 2890 1 5654
2 2891 1 5654
2 2892 1 5654
2 2893 1 5654
2 2894 1 5654
2 2895 1 5654
2 2896 1 5654
2 2897 1 5654
2 2898 1 5670
2 2899 1 5670
2 2900 1 5670
2 2901 1 5670
2 2902 1 5670
2 2903 1 5670
2 2904 1 5670
2 2905 1 5670
2 2906 1 5670
2 2907 1 5670
2 2908 1 5670
2 2909 1 5670
2 2910 1 5683
2 2911 1 5683
2 2912 1 5683
2 2938 1 5683
2 2939 1 5683
2 2940 1 5683
2 2941 1 5690
2 2942 1 5690
2 2943 1 5690
2 2944 1 5690
2 2945 1 5690
2 2946 1 5690
2 2947 1 5697
2 2948 1 5697
2 2949 1 5697
2 2950 1 5697
2 2951 1 5697
2 2952 1 5697
2 2953 1 5697
2 2954 1 5697
2 2955 1 5697
2 2956 1 5707
2 2957 1 5707
2 2958 1 5707
2 2959 1 5707
2 2960 1 5707
2 2961 1 5707
2 2962 1 5707
2 2963 1 5707
2 2964 1 5707
2 2965 1 5707
2 2966 1 5718
2 2967 1 5718
2 2968 1 5718
2 2969 1 5718
2 2970 1 5718
2 2971 1 5718
2 2972 1 5718
2 2973 1 5718
2 2974 1 5718
2 2975 1 5728
2 2976 1 5728
2 2977 1 5728
2 2978 1 5728
2 2979 1 5728
2 2980 1 5728
2 2981 1 5736
2 2982 1 5736
2 2983 1 5736
2 2984 1 5740
2 2985 1 5740
2 2986 1 5740
2 2987 1 5744
2 2989 1 5744
2 2990 1 5747
2 2991 1 5747
2 2992 1 5747
2 2993 1 5751
2 2994 1 5751
2 2995 1 5751
2 2996 1 5755
2 2997 1 5755
2 2998 1 5758
2 2999 1 5758
2 3000 1 5758
2 3001 1 5762
2 3002 1 5762
2 3003 1 5762
2 3004 1 5766
2 3010 1 5766
2 3011 1 5771
2 3012 1 5771
2 3013 1 5771
2 3014 1 5771
2 3015 1 5771
2 3016 1 5771
2 3017 1 5778
2 3018 1 5778
2 3019 1 5778
2 3030 1 5778
2 3031 1 5778
2 3042 1 5778
2 3043 1 5778
2 3044 1 5778
2 3045 1 5778
2 3046 1 5778
2 3047 1 5789
2 3048 1 5789
2 3049 1 5789
2 3050 1 5789
2 3051 1 5789
2 3052 1 5789
2 3053 1 5789
2 3054 1 5789
2 3055 1 5789
2 3056 1 5799
2 3057 1 5799
2 3058 1 5799
2 3059 1 5799
2 3060 1 5799
2 3062 1 5799
2 3063 1 5799
2 3065 1 5807
2 3066 1 5807
2 3068 1 5807
2 3069 1 5807
2 3071 1 5807
2 3072 1 5807
2 3074 1 5807
2 3075 1 5807
2 3076 1 5807
2 3077 1 5807
2 3078 1 5807
2 3079 1 5807
2 3081 1 5807
2 3082 1 5821
2 3083 1 5821
2 3084 1 5821
2 3085 1 5821
2 3086 1 5821
2 3087 1 5821
2 3088 1 5821
2 3089 1 5821
2 3090 1 5821
2 3091 1 5821
2 3092 1 5821
2 3093 1 5821
2 3094 1 5821
2 3095 1 5821
2 3098 1 5821
2 3099 1 5837
2 3100 1 5837
2 3102 1 5837
2 3103 1 5837
2 3104 1 5837
2 3105 1 5837
2 3106 1 5837
2 3108 1 5837
2 3109 1 5837
2 3110 1 5837
2 3111 1 5837
2 3112 1 5837
2 3113 1 5850
2 3115 1 5850
2 3116 1 5850
2 3117 1 5850
2 3118 1 5850
2 3119 1 5856
2 3120 1 5856
2 3121 1 5856
2 3123 1 5856
2 3124 1 5856
2 3125 1 5856
2 3127 1 5863
2 3128 1 5863
2 3129 1 5863
2 3132 1 5863
2 3133 1 5863
2 3138 1 5863
2 3139 1 5870
2 3141 1 5870
2 3142 1 5870
2 3143 1 5870
2 3145 1 5870
2 3146 1 5870
2 3147 1 5870
2 3148 1 5870
2 3150 1 5870
2 3151 1 5870
2 3152 1 5881
2 3153 1 5881
2 3154 1 5881
2 3156 1 5881
2 3157 1 5881
2 3158 1 5881
2 3160 1 5881
2 3161 1 5881
2 3162 1 5881
2 3163 1 5881
2 3164 1 5892
2 3165 1 5892
2 3166 1 5892
2 3170 1 5892
2 3171 1 5892
2 3172 1 5898
2 3174 1 5898
2 3175 1 5898
2 3176 1 5898
2 3177 1 5898
2 3179 1 5898
2 3180 1 5905
2 3181 1 5905
2 3182 1 5905
2 3183 1 5905
2 3186 1 5905
2 3187 1 5905
2 3188 1 5905
2 3190 1 5905
2 3191 1 5905
2 3192 1 5915
2 3193 1 5915
2 3194 1 5915
2 3196 1 5915
2 3197 1 5915
2 3198 1 5915
2 3199 1 5915
2 3200 1 5915
2 3201 1 5915
2 3203 1 5915
2 3204 1 5926
2 3205 1 5926
2 3206 1 5926
2 3207 1 5926
2 3208 1 5926
2 3209 1 5926
2 3212 1 5926
2 3213 1 5926
2 3214 1 5926
2 3216 1 5936
2 3217 1 5936
2 3218 1 5936
2 3219 1 5936
2 3220 1 5936
2 3222 1 5936
2 3223 1 5960
2 3224 1 5960
2 3225 1 5960
2 3226 1 5960
2 3227 1 5960
2 3230 1 5981
2 3231 1 5981
2 3233 1 5981
2 3234 1 5981
2 3235 1 5981
2 3237 1 5981
2 3238 1 5981
2 3239 1 5991
2 3240 1 5991
2 3242 1 5991
2 3243 1 5991
2 3244 1 5996
2 3245 1 5996
2 3246 1 5996
2 3248 1 6000
2 3249 1 6000
2 3250 1 6003
2 3252 1 6003
2 3253 1 6003
2 3254 1 6003
2 3256 1 6003
2 3257 1 6009
2 3258 1 6009
2 3260 1 6009
2 3261 1 6009
2 3262 1 6014
2 3264 1 6014
2 3265 1 6014
2 3266 1 6018
2 3268 1 6018
2 3269 1 6041
2 3270 1 6041
2 3271 1 6041
2 3272 1 6041
2 3274 1 6041
2 3275 1 6047
2 3276 1 6047
2 3277 1 6047
2 3278 1 6047
2 3279 1 6052
2 3280 1 6052
2 3282 1 6052
2 3283 1 6056
2 3284 1 6056
2 3285 1 6079
2 3286 1 6079
2 3288 1 6079
2 3289 1 6083
2 3290 1 6083
2 3291 1 6083
2 3292 1 6087
2 3294 1 6087
2 3295 1 6127
2 3296 1 6127
2 3297 1 6127
2 3298 1 6131
2 3300 1 6131
2 3301 1 6131
2 3302 1 6137
2 3304 1 6137
2 3305 1 6137
2 3306 1 6141
2 3308 1 6141
2 3309 1 6141
2 3310 1 6145
2 3312 1 6145
2 3313 1 6166
2 3314 1 6166
2 3316 1 6166
2 3317 1 6170
2 3318 1 6170
2 3319 1 6170
2 3320 1 6174
2 3321 1 6174
2 3323 1 6177
2 3324 1 6177
2 3325 1 6177
2 3326 1 6196
2 3327 1 6196
2 3329 1 6199
2 3330 1 6199
2 3331 1 6204
2 3332 1 6204
2 3333 1 6207
2 3335 1 6207
2 3336 1 6210
2 3337 1 6210
2 3338 1 6214
2 3339 1 6214
2 3341 1 6217
2 3342 1 6217
2 3344 1 6220
2 3345 1 6220
2 3346 1 6232
2 3347 1 6232
2 3348 1 6236
2 3350 1 6236
2 3351 1 6243
2 3352 1 6243
2 3353 1 6246
2 3354 1 6246
2 3356 1 6249
2 3357 1 6249
2 3358 1 6252
2 3359 1 6252
2 3360 1 6263
2 3376 1 6263
2 3377 1 6266
2 3378 1 6266
2 3382 1 6762
2 3383 1 6762
2 3385 1 6762
2 3386 1 6784
2 3387 1 6784
2 3388 1 6797
2 3389 1 6797
2 3391 1 6800
2 3392 1 6800
2 3393 1 6803
2 3394 1 6803
2 3395 1 6806
2 3396 1 6806
2 3397 1 6809
2 3399 1 6809
2 3400 1 6812
2 3401 1 6812
2 3402 1 6815
2 3403 1 6815
2 3405 1 6818
2 3406 1 6818
2 3407 1 6821
2 3408 1 6821
2 3409 1 6824
2 3411 1 6824
2 3412 1 6827
2 3413 1 6827
2 3414 1 6830
2 3415 1 6830
2 3417 1 6833
2 3418 1 6833
2 3419 1 6845
2 3421 1 6845
2 3422 1 6867
2 3423 1 6867
2 3425 1 6881
2 3426 1 6881
2 3427 1 6894
2 3429 1 6894
2 3430 1 6894
2 3431 1 6894
2 3433 1 6894
2 3434 1 6894
2 3435 1 6901
2 3437 1 6901
2 3438 1 6901
2 3439 1 6901
2 3441 1 6901
2 3442 1 6901
2 3443 1 6901
2 3445 1 6901
2 3446 1 6901
2 3447 1 6901
2 3449 1 6912
2 3450 1 6912
2 3451 1 6912
2 3455 1 6912
2 3456 1 6912
2 3457 1 6912
2 3459 1 6912
2 3460 1 6912
2 3461 1 6912
2 3463 1 6912
2 3464 1 6923
2 3465 1 6923
2 3467 1 6923
2 3468 1 6923
2 3469 1 6923
2 3471 1 6929
2 3472 1 6929
2 3473 1 6929
2 3475 1 6929
2 3476 1 6929
2 3477 1 6929
2 3479 1 6936
2 3480 1 6936
2 3481 1 6936
2 3483 1 6936
2 3484 1 6936
2 3485 1 6936
2 3488 1 6936
2 3489 1 6936
2 3491 1 6936
2 3492 1 6946
2 3494 1 6946
2 3495 1 6946
2 3497 1 6946
2 3498 1 6946
2 3500 1 6946
2 3501 1 6946
2 3503 1 6946
2 3504 1 6946
2 3505 1 6946
2 3506 1 6957
2 3508 1 6957
2 3509 1 6957
2 3511 1 6957
2 3512 1 6957
2 3513 1 6957
2 3514 1 6957
2 3516 1 6957
2 3517 1 6957
2 3519 1 6970
2 3520 1 6970
2 3522 1 6970
2 3523 1 6970
2 3525 1 6970
2 3526 1 6970
2 3528 1 6977
2 3529 1 6977
2 3531 1 6977
2 3532 1 6977
2 3533 1 6977
2 3534 1 6977
2 3536 1 6977
2 3537 1 6977
2 3538 1 6977
2 3540 1 6977
2 3541 1 6988
2 3543 1 6988
2 3544 1 6988
2 3546 1 6988
2 3547 1 6988
2 3549 1 6988
2 3550 1 6988
2 3554 1 6988
2 3555 1 6988
2 3556 1 6998
2 3558 1 6998
2 3559 1 6998
2 3561 1 6998
2 3562 1 6998
2 3564 1 6998
2 3565 1 6998
2 3567 1 7006
2 3568 1 7006
2 3572 1 7006
2 3573 1 7006
2 3575 1 7006
2 3576 1 7006
2 3578 1 7006
2 3579 1 7006
2 3581 1 7006
2 3582 1 7006
2 3584 1 7006
2 3585 1 7006
2 3587 1 7006
2 3588 1 7020
2 3590 1 7020
2 3591 1 7020
2 3593 1 7020
2 3594 1 7020
2 3596 1 7020
2 3597 1 7020
2 3599 1 7020
2 3600 1 7020
2 3602 1 7020
2 3603 1 7020
2 3605 1 7020
2 3606 1 7020
2 3608 1 7020
2 3609 1 7020
2 3611 1 7036
2 3612 1 7036
2 3614 1 7036
2 3615 1 7036
2 3617 1 7036
2 3618 1 7036
2 3620 1 7036
2 3621 1 7036
2 3623 1 7036
2 3624 1 7036
2 3626 1 7036
2 3627 1 7036
2 3629 1 7049
2 3630 1 7049
2 3632 1 7049
2 3633 1 7049
2 3635 1 7049
2 3636 1 7057
2 3638 1 7057
2 3639 1 7068
2 3641 1 7068
2 3642 1 7068
2 3644 1 7068
2 3645 1 7073
2 3647 1 7073
2 3648 1 7073
2 3650 1 7077
2 3651 1 7077
2 3653 1 7080
2 3654 1 7080
2 3656 1 7080
2 3657 1 7080
2 3659 1 7080
2 3660 1 7086
2 3662 1 7086
2 3663 1 7086
2 3665 1 7086
2 3666 1 7091
2 3668 1 7091
2 3669 1 7091
2 3671 1 7095
2 3672 1 7095
2 3674 1 7100
2 3675 1 7100
2 3677 1 7107
2 3678 1 7107
2 3680 1 7107
2 3681 1 7107
2 3683 1 7107
2 3684 1 7107
2 3686 1 7114
2 3687 1 7114
2 3689 1 7114
2 3690 1 7114
2 3692 1 7114
2 3693 1 7114
2 3695 1 7114
2 3696 1 7114
2 3698 1 7114
2 3699 1 7114
2 3701 1 7125
2 3702 1 7125
2 3704 1 7125
2 3705 1 7125
2 3707 1 7125
2 3708 1 7125
2 3710 1 7125
2 3711 1 7125
2 3713 1 7125
2 3714 1 7125
2 3716 1 7136
2 3717 1 7136
2 3719 1 7136
2 3720 1 7136
2 3722 1 7136
2 3723 1 7142
2 3725 1 7142
2 3726 1 7142
2 3728 1 7142
2 3729 1 7142
2 3731 1 7142
2 3732 1 7149
2 3734 1 7149
2 3735 1 7149
2 3737 1 7149
2 3738 1 7149
2 3740 1 7149
2 3741 1 7149
2 3743 1 7149
2 3744 1 7149
2 3746 1 7159
2 3747 1 7159
2 3749 1 7159
2 3750 1 7159
2 3752 1 7159
2 3753 1 7159
2 3755 1 7159
2 3756 1 7159
2 3758 1 7159
2 3759 1 7159
2 3761 1 7170
2 3762 1 7170
2 3764 1 7170
2 3765 1 7170
2 3767 1 7170
2 3768 1 7170
2 3770 1 7170
2 3771 1 7170
2 3773 1 7170
2 3774 1 7180
2 3776 1 7180
2 3777 1 7180
2 3779 1 7180
2 3780 1 7180
2 3784 1 7180
2 3785 1 7188
2 3787 1 7188
2 3788 1 7191
2 3790 1 7191
2 3791 1 7194
2 3793 1 7194
2 3794 1 7194
2 3796 1 7198
2 3797 1 7198
2 3799 1 7198
2 3800 1 7202
2 3802 1 7202
2 3803 1 7205
2 3805 1 7205
2 3806 1 7205
2 3808 1 7209
2 3809 1 7209
2 3811 1 7209
2 3812 1 7213
2 3814 1 7213
2 3815 1 7216
2 3817 1 7216
2 3818 1 7219
2 3820 1 7219
2 3821 1 7222
2 3823 1 7222
2 3824 1 7222
2 3826 1 7222
2 3827 1 7222
2 3829 1 7222
2 3830 1 7229
2 3832 1 7229
2 3833 1 7229
2 3835 1 7229
2 3836 1 7229
2 3838 1 7229
2 3839 1 7229
2 3841 1 7229
2 3842 1 7229
2 3844 1 7229
2 3845 1 7240
2 3847 1 7240
2 3848 1 7240
2 3850 1 7240
2 3851 1 7240
2 3853 1 7240
2 3854 1 7240
2 3856 1 7240
2 3857 1 7240
2 3859 1 7250
2 3860 1 7250
2 3862 1 7250
2 3863 1 7250
2 3865 1 7250
2 3866 1 7250
2 3868 1 7250
2 3869 1 7258
2 3871 1 7258
2 3872 1 7258
2 3874 1 7258
2 3875 1 7258
2 3877 1 7258
2 3878 1 7258
2 3880 1 7258
2 3881 1 7258
2 3883 1 7258
2 3884 1 7258
2 3886 1 7258
2 3887 1 7258
2 3889 1 7272
2 3890 1 7272
2 3892 1 7272
2 3893 1 7272
2 3894 1 7272
2 3895 1 7272
2 3896 1 7272
2 3897 1 7272
2 3898 1 7272
2 3899 1 7272
2 3900 1 7272
2 3901 1 7272
2 3902 1 7272
2 3903 1 7272
2 3904 1 7272
2 3905 1 7288
2 3906 1 7288
2 3907 1 7288
2 3908 1 7288
2 3909 1 7288
2 3910 1 7288
2 3911 1 7288
2 3912 1 7288
2 3913 1 7288
2 3914 1 7288
2 3915 1 7288
2 3916 1 7288
2 3917 1 7301
2 3918 1 7301
2 3919 1 7301
2 3920 1 7301
2 3921 1 7301
2 3922 1 7307
2 3923 1 7307
2 3924 1 7307
2 3925 1 7307
2 3926 1 7307
2 3927 1 7307
2 3928 1 7314
2 3929 1 7314
2 3930 1 7314
2 3931 1 7318
2 3932 1 7318
2 3933 1 7318
2 3934 1 7322
2 3935 1 7322
2 3936 1 7325
2 3937 1 7325
2 3938 1 7328
2 3939 1 7328
2 3940 1 7331
2 3941 1 7331
2 3942 1 7334
2 3943 1 7334
2 3944 1 7337
2 3945 1 7337
2 3946 1 7340
2 3947 1 7340
2 3948 1 7343
2 3949 1 7343
2 3950 1 7346
2 3951 1 7346
2 3952 1 7346
2 3957 1 7346
2 3959 1 7351
2 3960 1 7351
2 3961 1 7351
2 3962 1 7355
2 3963 1 7355
2 3965 1 7358
2 3966 1 7358
2 3967 1 7358
2 3968 1 7358
2 3969 1 7358
2 3970 1 7364
2 3971 1 7364
2 3972 1 7364
2 3973 1 7364
2 3974 1 7369
2 3975 1 7369
2 3976 1 7369
2 3977 1 7373
2 3978 1 7373
2 3979 1 7378
2 3980 1 7378
2 3981 1 7381
2 3982 1 7381
2 3983 1 7384
2 3984 1 7384
2 3985 1 7387
2 3986 1 7387
2 3987 1 7387
2 3988 1 7391
2 3989 1 7391
2 3990 1 7394
2 3991 1 7394
2 3992 1 7394
2 3993 1 7398
2 3994 1 7398
2 3995 1 7398
2 3996 1 7402
2 3997 1 7402
2 3998 1 7405
2 3999 1 7405
2 4000 1 7408
2 4001 1 7408
2 4002 1 7411
2 4003 1 7411
2 4004 1 7414
2 4005 1 7414
2 4006 1 7417
2 4007 1 7417
2 4008 1 7420
2 4009 1 7420
2 4010 1 7423
2 4011 1 7423
2 4012 1 7426
2 4013 1 7426
2 4014 1 7429
2 4015 1 7429
2 4016 1 7432
2 4017 1 7432
2 4018 1 7435
2 4019 1 7435
2 4020 1 7438
2 4021 1 7438
2 4022 1 7441
2 4023 1 7441
2 4024 1 7444
2 4025 1 7444
2 4026 1 7447
2 4027 1 7447
2 4028 1 7450
2 4029 1 7450
2 4030 1 7453
2 4031 1 7453
2 4032 1 7456
2 4033 1 7456
2 4034 1 7459
2 4035 1 7459
2 4036 1 7462
2 4037 1 7462
2 4038 1 7465
2 4039 1 7465
2 4040 1 7468
2 4041 1 7468
2 4042 1 7471
2 4043 1 7471
2 4044 1 7474
2 4045 1 7474
2 4046 1 7479
2 4047 1 7479
2 4048 1 7482
2 4049 1 7482
2 4050 1 7485
2 4051 1 7485
2 4052 1 7488
2 4053 1 7488
2 4054 1 7491
2 4055 1 7491
2 4056 1 7494
2 4057 1 7494
2 4058 1 7497
2 4059 1 7497
2 4060 1 7500
2 4061 1 7500
2 4062 1 7503
2 4063 1 7503
2 4064 1 7506
2 4065 1 7506
2 4066 1 7509
2 4067 1 7509
2 4068 1 7512
2 4069 1 7512
2 4070 1 7515
2 4071 1 7515
2 4072 1 7518
2 4073 1 7518
2 4074 1 7521
2 4075 1 7521
2 4076 1 7524
2 4077 1 7524
2 4078 1 7527
2 4079 1 7527
2 4080 1 7530
2 4081 1 7530
2 4082 1 7533
2 4083 1 7533
2 4084 1 7536
2 4085 1 7536
2 4086 1 7539
2 4087 1 7539
2 4088 1 7542
2 4089 1 7542
2 4090 1 7545
2 4091 1 7545
2 4092 1 7548
2 4093 1 7548
2 4094 1 7553
2 4095 1 7553
2 4096 1 7560
2 4097 1 7560
2 4098 1 7563
2 4099 1 7563
2 4100 1 7566
2 4101 1 7566
2 4102 1 7569
2 4103 1 7569
2 4104 1 7574
2 4105 1 7574
2 4106 1 7577
2 4107 1 7577
2 4108 1 7582
2 4109 1 7582
2 4110 1 7585
2 4111 1 7585
2 4112 1 7588
2 4113 1 7588
2 4114 1 7591
2 4115 1 7591
2 4116 1 7609
2 4117 1 7609
2 4118 1 7609
2 4119 1 7613
2 4120 1 7613
2 4121 1 7620
2 4122 1 7620
2 4123 1 7650
2 4124 1 7650
2 4125 1 7655
2 4126 1 7655
2 4127 1 7655
2 4128 1 7659
2 4129 1 7659
2 4130 1 7671
2 4131 1 7671
2 4132 1 7852
2 4133 1 7852
2 4134 1 8114
2 4135 1 8114
2 4136 1 8117
2 4137 1 8117
2 4138 1 8131
2 4139 1 8131
2 4140 1 8134
2 4141 1 8134
2 4142 1 8146
2 4143 1 8146
2 4144 1 8156
2 4145 1 8156
2 4146 1 8166
2 4147 1 8166
2 4148 1 8169
2 4149 1 8169
2 4150 1 8183
2 4151 1 8183
2 4152 1 8186
2 4153 1 8186
2 4154 1 8196
2 4155 1 8196
2 4156 1 8200
2 4157 1 8200
2 4158 1 8204
2 4159 1 8204
2 4160 1 8208
2 4161 1 8208
2 4162 1 8262
2 4163 1 8262
2 4164 1 8262
2 4165 1 8262
2 4166 1 8269
2 4167 1 8269
2 4168 1 8269
2 4169 1 8269
2 4170 1 8298
2 4171 1 8298
2 4172 1 8298
2 4173 1 8298
2 4174 1 8298
2 4175 1 8298
2 4176 1 8307
2 4177 1 8307
2 4178 1 8307
2 4179 1 8307
2 4180 1 8307
2 4181 1 8307
2 4182 1 8326
2 4183 1 8326
2 4184 1 8326
2 4185 1 8326
2 4186 1 8326
2 4187 1 8326
2 4188 1 8333
2 4189 1 8333
2 4190 1 8333
2 4191 1 8358
2 4192 1 8358
2 4194 1 8358
2 4195 1 8358
2 4196 1 8358
2 4197 1 8358
2 4198 1 8365
2 4199 1 8365
2 4200 1 8365
2 4201 1 8394
2 4202 1 8394
2 4203 1 8394
2 4204 1 8394
2 4205 1 8394
2 4206 1 8394
2 4207 1 8394
2 4208 1 8394
2 4209 1 8394
2 4210 1 8405
2 4211 1 8405
2 4212 1 8405
2 4213 1 8412
2 4214 1 8412
2 4215 1 8421
2 4216 1 8421
2 4217 1 8421
2 4218 1 8421
2 4219 1 8421
2 4220 1 8421
2 4221 1 8421
2 4222 1 8421
2 4223 1 8430
2 4224 1 8430
2 4225 1 8444
2 4226 1 8444
2 4227 1 8457
2 4228 1 8457
2 4229 1 8460
2 4230 1 8460
2 4231 1 8463
2 4232 1 8463
2 4233 1 8466
2 4234 1 8466
2 4235 1 8471
2 4236 1 8471
2 4237 1 8474
2 4238 1 8474
2 4239 1 8477
2 4240 1 8477
2 4241 1 8480
2 4242 1 8480
2 4243 1 8485
2 4244 1 8485
2 4245 1 8497
2 4246 1 8497
2 4247 1 8519
2 4248 1 8519
2 4249 1 8522
2 4250 1 8522
2 4251 1 8525
2 4252 1 8525
2 4253 1 8528
2 4254 1 8528
2 4255 1 8531
2 4256 1 8531
2 4257 1 8534
2 4258 1 8534
2 4259 1 8541
2 4260 1 8541
2 4261 1 8541
2 4262 1 8548
2 4263 1 8548
2 4264 1 8555
2 4265 1 8555
2 4266 1 8558
2 4267 1 8558
2 4268 1 8561
2 4269 1 8561
2 4270 1 8566
2 4271 1 8566
2 4272 1 8569
2 4273 1 8569
2 4274 1 8572
2 4275 1 8572
2 4276 1 8575
2 4277 1 8575
2 4278 1 8580
2 4279 1 8580
2 4280 1 8583
2 4281 1 8583
2 4282 1 8586
2 4283 1 8586
2 4284 1 8589
2 4285 1 8589
2 4286 1 8592
2 4287 1 8592
2 4288 1 8595
2 4289 1 8595
2 4290 1 8598
2 4291 1 8598
2 4292 1 8601
2 4293 1 8601
2 4294 1 8604
2 4295 1 8604
2 4296 1 8627
2 4297 1 8627
2 4298 1 8660
2 4299 1 8660
2 4300 1 8663
2 4301 1 8663
2 4302 1 8666
2 4304 1 8666
2 4305 1 8669
2 4306 1 8669
2 4307 1 8672
2 4309 1 8672
2 4310 1 8675
2 4311 1 8675
2 4312 1 8678
2 4314 1 8678
2 4315 1 8681
2 4316 1 8681
2 4317 1 8684
2 4318 1 8684
2 4319 1 8687
2 4320 1 8687
2 4321 1 8690
2 4322 1 8690
2 4323 1 8693
2 4324 1 8693
2 4325 1 8696
2 4328 1 8696
2 4329 1 8699
2 4330 1 8699
2 4331 1 8702
2 4332 1 8702
2 4335 1 8705
2 4336 1 8705
2 4337 1 8708
2 4338 1 8708
2 4339 1 8711
2 4340 1 8711
2 4341 1 8714
2 4342 1 8714
2 4343 1 8718
2 4344 1 8718
2 4345 1 8721
2 4346 1 8721
2 4347 1 8724
2 4348 1 8724
2 4349 1 8727
2 4350 1 8727
2 4351 1 8730
2 4352 1 8730
2 4353 1 8735
2 4354 1 8735
2 4355 1 8738
2 4356 1 8738
2 4357 1 8741
2 4358 1 8741
2 4359 1 8744
2 4360 1 8744
2 4361 1 8747
2 4362 1 8747
2 4363 1 8750
2 4364 1 8750
2 4365 1 8757
2 4366 1 8757
2 4367 1 8760
2 4368 1 8760
2 4369 1 8763
2 4370 1 8763
2 4371 1 8766
2 4372 1 8766
2 4373 1 8769
2 4374 1 8769
2 4375 1 8772
2 4376 1 8772
2 4377 1 8775
2 4378 1 8775
2 4379 1 8778
2 4380 1 8778
2 4381 1 8781
2 4382 1 8781
2 4383 1 8784
2 4384 1 8784
2 4385 1 8787
2 4386 1 8787
2 4387 1 8790
2 4388 1 8790
2 4389 1 8793
2 4390 1 8793
2 4391 1 8796
2 4392 1 8796
2 4393 1 8799
2 4394 1 8799
2 4395 1 8802
2 4396 1 8802
2 4397 1 8805
2 4398 1 8805
2 4399 1 8808
2 4400 1 8808
2 4401 1 8811
2 4402 1 8811
2 4403 1 8857
2 4404 1 8857
2 4405 1 8857
2 4406 1 8871
2 4407 1 8871
2 4408 1 8898
2 4409 1 8898
2 4410 1 8898
2 4413 1 8902
2 4414 1 8902
2 4415 1 8920
2 4416 1 8920
2 4417 1 8920
2 4418 1 8924
2 4419 1 8924
2 4420 1 8927
2 4421 1 8927
2 4422 1 8927
2 4423 1 8931
2 4424 1 8931
2 4425 1 8943
2 4426 1 8943
2 4427 1 8943
2 4428 1 8950
2 4429 1 8950
2 4430 1 8950
2 4431 1 8956
2 4432 1 8956
2 4433 1 8966
2 4434 1 8966
2 4435 1 8996
2 4436 1 8996
2 4437 1 9001
2 4438 1 9001
2 4439 1 9001
2 4440 1 9005
2 4441 1 9005
2 4442 1 9029
2 4443 1 9029
2 4444 1 9029
2 4445 1 9035
2 4446 1 9035
2 4447 1 9068
2 4448 1 9068
2 4449 1 9074
2 4450 1 9074
2 4451 1 9079
2 4452 1 9079
2 4453 1 9083
2 4454 1 9083
2 4455 1 9089
2 4456 1 9089
2 4457 1 9095
2 4458 1 9095
2 4459 1 9099
2 4460 1 9099
2 4461 1 9103
2 4462 1 9103
2 4546 1 9107
2 4547 1 9107
2 4548 1 9111
2 4550 1 9111
2 4551 1 9117
2 4552 1 9117
2 4553 1 9127
2 4554 1 9127
2 4556 1 9146
2 4557 1 9146
2 4558 1 9149
2 4559 1 9149
2 4560 1 9161
2 4561 1 9161
2 4564 1 9165
2 4565 1 9165
2 4567 1 9169
2 4568 1 9169
2 4569 1 9173
2 4571 1 9173
2 4572 1 9183
2 4573 1 9183
2 4574 1 9193
2 4578 1 9193
2 4579 1 9203
2 4580 1 9203
2 4582 1 9206
2 4583 1 9206
2 4584 1 9220
2 4585 1 9220
2 4587 1 9223
2 4588 1 9223
2 4589 1 9265
2 4590 1 9265
2 4591 1 9268
2 4594 1 9268
2 4595 1 9280
2 4596 1 9280
2 4598 1 9307
2 4599 1 9307
2 4600 1 9307
2 4601 1 9332
2 4602 1 9332
2 4604 1 9332
2 4605 1 9332
2 4606 1 9332
2 4607 1 9332
2 4608 1 9339
2 4609 1 9339
2 4654 1 9344
2 4655 1 9344
2 4658 1 9344
2 4659 1 9344
2 4660 1 9344
2 4662 1 9344
2 4663 1 9385
2 4664 1 9385
2 4665 1 9385
2 4666 1 9385
2 4668 1 9385
2 4669 1 9385
2 4670 1 9408
2 4671 1 9408
2 4672 1 9408
2 4673 1 9423
2 4676 1 9423
2 4677 1 9426
2 4679 1 9426
2 4680 1 9429
2 4681 1 9429
2 4683 1 9462
2 4684 1 9462
2 4685 1 9473
2 4686 1 9473
2 4688 1 9478
2 4689 1 9478
2 4690 1 9485
2 4691 1 9485
2 4692 1 9488
2 4703 1 9488
2 4704 1 9517
2 4705 1 9517
2 4707 1 9520
2 4708 1 9520
2 4709 1 9543
2 4710 1 9543
2 4712 1 9551
2 4713 1 9551
2 4714 1 9575
2 4715 1 9575
2 4716 1 9575
2 4719 1 9608
2 4720 1 9608
2 4721 1 9626
2 4723 1 9626
2 4724 1 9629
2 4725 1 9629
2 4726 1 9632
2 4727 1 9632
2 4729 1 9635
2 4730 1 9635
2 4731 1 9642
2 4732 1 9642
2 4733 1 9646
2 4734 1 9646
2 4736 1 9650
2 4737 1 9650
2 4738 1 9653
2 4739 1 9653
2 4740 1 9656
2 4741 1 9656
2 4742 1 9663
2 4770 1 9663
2 4771 1 9667
2 4772 1 9667
2 4773 1 9671
2 4774 1 9671
2 4785 1 9675
2 4786 1 9675
2 4787 1 9679
2 4788 1 9679
2 4791 1 9682
2 4792 1 9682
2 4797 1 9685
2 4798 1 9685
2 4804 1 9692
2 4805 1 9692
2 4807 1 9698
2 4808 1 9698
2 4811 1 9702
2 4812 1 9702
2 4815 1 9707
2 4816 1 9707
2 4818 1 9711
2 4819 1 9711
2 4821 1 9717
2 4822 1 9717
2 4824 1 9723
2 4825 1 9723
2 4827 1 9727
2 4828 1 9727
2 4830 1 9754
2 4831 1 9754
2 4833 1 9754
2 4834 1 9758
2 4836 1 9758
2 4837 1 9758
2 4839 1 9775
2 4840 1 9775
2 4842 1 9775
2 4843 1 9779
2 4845 1 9779
2 4846 1 9779
2 4848 1 9786
2 4849 1 9786
2 4851 1 9786
2 4852 1 9791
2 4854 1 9791
2 4855 1 9791
2 4857 1 9809
2 4858 1 9809
2 4860 1 9809
2 4861 1 9817
2 4863 1 9817
2 4864 1 9820
2 4866 1 9820
2 4867 1 9820
2 4869 1 9925
2 4870 1 9925
2 4872 1 9925
2 4873 1 9925
2 4875 1 9925
2 4876 1 9925
2 4878 1 9932
2 4879 1 9932
2 4881 1 9935
2 4882 1 9935
2 4884 1 9949
2 4885 1 9949
2 4887 1 9961
2 4888 1 9961
2 4890 1 9964
2 4891 1 9964
2 4893 1 9979
2 4894 1 9979
2 4896 1 9983
2 4897 1 9983
2 4899 1 9986
2 4900 1 9986
2 4902 1 9989
2 4903 1 9989
2 4905 1 9992
2 4906 1 9992
2 4908 1 9999
2 4909 1 9999
2 4911 1 10003
2 4912 1 10003
2 4914 1 10007
2 4915 1 10007
2 4917 1 10010
2 4918 1 10010
2 4920 1 10070
2 4921 1 10070
2 4923 1 10073
2 4924 1 10073
2 4926 1 10116
2 4927 1 10116
2 4929 1 10119
2 4930 1 10119
2 4932 1 10119
2 4933 1 10119
2 4935 1 10124
2 4936 1 10124
2 4938 1 10124
2 4939 1 10124
2 4941 1 10124
2 4942 1 10141
2 4944 1 10141
2 4945 1 10141
2 4947 1 10141
2 4948 1 10141
2 4950 1 10141
2 4951 1 10148
2 4953 1 10148
2 4954 1 10148
2 4956 1 10148
2 4957 1 10148
2 4959 1 10148
2 4960 1 10170
2 4962 1 10170
2 4963 1 10173
2 4965 1 10173
2 4966 1 10180
2 4968 1 10180
2 4969 1 10183
2 4971 1 10183
2 4972 1 10186
2 4974 1 10186
2 4975 1 10189
2 4977 1 10189
2 4978 1 10192
2 4980 1 10192
2 4981 1 10197
2 4983 1 10197
2 4984 1 10200
2 4986 1 10200
2 4987 1 10273
2 4989 1 10273
2 4990 1 10273
2 4992 1 10273
2 4993 1 10283
2 4995 1 10283
2 4996 1 10283
2 4998 1 10296
2 4999 1 10296
2 5001 1 10301
2 5002 1 10301
2 5004 1 10301
2 5005 1 10301
2 5007 1 10308
2 5008 1 10308
2 5010 1 10311
2 5011 1 10311
2 5013 1 10318
2 5014 1 10318
2 5016 1 10321
2 5017 1 10321
2 5019 1 10334
2 5020 1 10334
2 5022 1 10341
2 5023 1 10341
2 5025 1 10344
2 5026 1 10344
2 5028 1 10354
2 5029 1 10354
2 5031 1 10357
2 5032 1 10357
2 5034 1 10360
2 5035 1 10360
2 5037 1 10367
2 5038 1 10367
2 5040 1 10367
2 5041 1 10367
2 5043 1 10375
2 5044 1 10375
2 5050 1 10375
2 5051 1 10375
2 5053 1 10375
2 5054 1 10381
2 5056 1 10381
2 5057 1 10381
2 5059 1 10381
2 5060 1 10381
2 5062 1 10381
2 5063 1 10388
2 5069 1 10388
2 5070 1 10391
2 5072 1 10391
2 5073 1 10399
2 5075 1 10399
2 5076 1 10402
2 5078 1 10402
2 5079 1 10406
2 5081 1 10406
2 5082 1 10409
2 5084 1 10409
2 5085 1 10412
2 5087 1 10412
2 5088 1 10415
2 5090 1 10415
2 5091 1 10419
2 5093 1 10419
2 5094 1 10422
2 5096 1 10422
2 5097 1 10425
2 5099 1 10425
2 5100 1 10428
2 5102 1 10428
2 5103 1 10479
2 5105 1 10479
2 5106 1 10479
2 5108 1 10497
2 5109 1 10497
2 5115 1 10497
2 5116 1 10509
2 5118 1 10509
2 5119 1 10512
2 5121 1 10512
2 5122 1 10519
2 5124 1 10519
2 5125 1 10522
2 5127 1 10522
2 5128 1 10525
2 5130 1 10525
2 5131 1 10528
2 5133 1 10528
2 5134 1 10531
2 5136 1 10531
2 5137 1 10536
2 5139 1 10536
2 5140 1 10539
2 5142 1 10539
2 5143 1 10583
2 5145 1 10583
2 5146 1 10583
2 5148 1 10589
2 5149 1 10589
2 5151 1 10589
2 5152 1 10589
2 5154 1 10602
2 5155 1 10602
2 5157 1 10652
2 5158 1 10652
2 5160 1 10652
2 5161 1 10652
2 5163 1 10652
2 5164 1 10659
2 5194 1 10659
2 5195 1 10662
2 5214 1 10662
2 5215 1 10665
2 5216 1 10665
2 5217 1 10668
2 5218 1 10668
2 5219 1 10675
2 5220 1 10675
2 5221 1 10678
2 5222 1 10678
2 5223 1 10691
2 5224 1 10691
2 5225 1 10698
2 5226 1 10698
2 5227 1 10701
2 5228 1 10701
2 5229 1 10739
2 5230 1 10739
2 5231 1 10778
2 5232 1 10778
2 5233 1 10781
2 5234 1 10781
2 5235 1 10784
2 5236 1 10784
2 5237 1 10784
2 5238 1 10784
2 5239 1 10789
2 5240 1 10789
2 5241 1 10792
2 5242 1 10792
2 5243 1 10800
2 5244 1 10800
2 5245 1 10803
2 5246 1 10803
2 5247 1 10806
2 5248 1 10806
2 5249 1 10809
2 5250 1 10809
2 5251 1 10812
2 5252 1 10812
2 5253 1 10817
2 5254 1 10817
2 5255 1 10820
2 5256 1 10820
2 5257 1 10876
2 5258 1 10876
2 5259 1 10879
2 5260 1 10879
2 5261 1 10892
2 5262 1 10892
2 5263 1 10899
2 5264 1 10899
2 5265 1 10902
2 5266 1 10902
2 5267 1 10928
2 5268 1 10928
2 5269 1 10931
2 5270 1 10931
2 5271 1 10938
2 5272 1 10938
2 5273 1 10941
2 5274 1 10941
2 5275 1 10944
2 5276 1 10944
2 5277 1 10947
2 5278 1 10947
2 5279 1 10950
2 5280 1 10950
2 5281 1 10955
2 5282 1 10955
2 5301 1 10958
2 5302 1 10958
2 5303 1 10992
2 5304 1 10992
2 5305 1 10995
2 5306 1 10995
2 5307 1 11008
2 5308 1 11008
2 5309 1 11015
2 5310 1 11015
2 5311 1 11018
2 5312 1 11018
2 5313 1 11044
2 5325 1 11044
2 5326 1 11047
2 5327 1 11047
2 5328 1 11050
2 5329 1 11050
2 5330 1 11053
2 5331 1 11053
2 5332 1 11056
2 5333 1 11056
2 5334 1 11059
2 5335 1 11059
2 5336 1 11062
2 5337 1 11062
2 5338 1 11067
2 5339 1 11067
2 5340 1 11070
2 5341 1 11070
2 5342 1 11100
2 5343 1 11100
2 5344 1 11103
2 5345 1 11103
2 5346 1 11124
2 5347 1 11124
2 5348 1 11127
2 5349 1 11127
2 5350 1 11130
2 5351 1 11130
2 5352 1 11156
2 5353 1 11156
2 5354 1 11159
2 5355 1 11159
2 5356 1 11162
2 5357 1 11162
2 5358 1 11165
2 5359 1 11165
2 5360 1 11168
2 5361 1 11168
2 5362 1 11171
2 5368 1 11171
2 5369 1 11174
2 5370 1 11174
2 5371 1 11177
2 5372 1 11177
2 5373 1 11180
2 5374 1 11180
2 5375 1 11205
2 5376 1 11205
2 5377 1 11233
2 5378 1 11233
2 5379 1 11236
2 5380 1 11236
2 5381 1 11239
2 5382 1 11239
2 5383 1 11252
2 5384 1 11252
2 5385 1 11257
2 5386 1 11257
2 5387 1 11272
2 5388 1 11272
2 5389 1 11299
2 5390 1 11299
2 5391 1 11302
2 5392 1 11302
2 5393 1 11317
2 5394 1 11317
2 5395 1 11323
2 5396 1 11323
