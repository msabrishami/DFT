1 1 0 1 0
1 2 0 1 0
1 3 0 1 0
1 4 0 1 0
1 5 0 1 0
1 6 0 1 0
1 7 0 1 0
1 8 0 2 0
1 11 0 2 0
1 14 0 1 0
1 15 0 1 0
1 16 0 2 0
1 19 0 1 0
1 20 0 1 0
1 21 0 1 0
1 22 0 1 0
1 23 0 1 0
1 24 0 1 0
1 25 0 1 0
1 26 0 1 0
1 27 0 1 0
1 28 0 1 0
1 29 0 2 0
1 32 0 1 0
1 33 0 1 0
1 34 0 1 0
1 35 0 1 0
1 36 0 1 0
1 37 0 2 0
1 40 0 2 0
1 43 0 1 0
1 44 0 2 0
1 47 0 1 0
1 48 0 1 0
1 49 0 1 0
1 50 0 1 0
1 51 0 1 0
1 52 0 1 0
1 53 0 1 0
1 54 0 1 0
1 55 0 1 0
1 56 0 1 0
1 57 0 2 0
1 60 0 1 0
1 61 0 1 0
1 62 0 1 0
1 63 0 1 0
1 64 0 1 0
1 65 0 1 0
1 66 0 1 0
1 67 0 1 0
1 68 0 1 0
1 69 0 2 0
1 72 0 1 0
1 73 0 1 0
1 74 0 1 0
1 75 0 1 0
1 76 0 1 0
1 77 0 1 0
1 78 0 1 0
1 79 0 1 0
1 80 0 1 0
1 81 0 1 0
1 82 0 2 0
1 85 0 1 0
1 86 0 1 0
1 87 0 1 0
1 88 0 1 0
1 89 0 1 0
1 90 0 1 0
1 91 0 1 0
1 92 0 1 0
1 93 0 1 0
1 94 0 1 0
1 95 0 1 0
1 96 0 2 0
1 99 0 1 0
1 100 0 1 0
1 101 0 1 0
1 102 0 1 0
1 103 0 1 0
1 104 0 1 0
1 105 0 1 0
1 106 0 1 0
1 107 0 1 0
1 108 0 2 0
1 111 0 1 0
1 112 0 1 0
1 113 0 1 0
1 114 0 1 0
1 115 0 1 0
1 116 0 1 0
1 117 0 1 0
1 118 0 1 0
1 119 0 1 0
1 120 0 2 0
1 123 0 1 0
1 124 0 1 0
1 125 0 1 0
1 126 0 1 0
1 127 0 1 0
1 128 0 1 0
1 129 0 1 0
1 130 0 1 0
1 131 0 1 0
1 132 0 2 0
1 135 0 1 0
1 136 0 1 0
1 137 0 1 0
1 138 0 1 0
1 139 0 1 0
1 140 0 1 0
1 141 0 1 0
1 142 0 1 0
3 143 0 0 0 
3 144 0 0 0 
3 145 0 0 0 
3 146 0 0 0 
3 147 0 0 0 
3 148 0 0 0 
3 149 0 0 0 
3 150 0 0 0 
3 151 0 0 0 
3 152 0 0 0 
3 153 0 0 0 
3 154 0 0 0 
3 155 0 0 0 
3 156 0 0 0 
3 157 0 0 0 
3 158 0 0 0 
3 159 0 0 0 
3 160 0 0 0 
3 161 0 0 0 
3 162 0 0 0 
3 163 0 0 0 
3 164 0 0 0 
3 165 0 0 0 
3 166 0 0 0 
3 167 0 0 0 
3 168 0 0 0 
3 169 0 0 0 
3 170 0 0 0 
3 171 0 0 0 
3 172 0 0 0 
3 173 0 0 0 
3 174 0 0 0 
3 175 0 0 0 
3 176 0 0 0 
3 177 0 0 0 
3 178 0 0 0 
3 179 0 0 0 
3 180 0 0 0 
3 181 0 0 0 
3 182 0 0 0 
3 183 0 0 0 
3 184 0 0 0 
3 185 0 0 0 
3 186 0 0 0 
3 187 0 0 0 
3 188 0 0 0 
3 189 0 0 0 
3 190 0 0 0 
3 191 0 0 0 
3 192 0 0 0 
3 193 0 0 0 
3 194 0 0 0 
3 195 0 0 0 
3 196 0 0 0 
3 197 0 0 0 
3 198 0 0 0 
3 199 0 0 0 
3 200 0 0 0 
3 201 0 0 0 
3 202 0 0 0 
3 203 0 0 0 
3 204 0 0 0 
3 205 0 0 0 
3 206 0 0 0 
3 207 0 0 0 
3 208 0 0 0 
3 209 0 0 0 
3 210 0 0 0 
3 211 0 0 0 
3 212 0 0 0 
3 213 0 0 0 
3 214 0 0 0 
3 215 0 0 0 
3 216 0 0 0 
3 217 0 0 0 
3 218 0 0 0 
1 219 0 4 0
1 224 0 2 0
1 227 0 2 0
1 230 0 1 0
1 231 0 2 0
1 234 0 2 0
1 237 0 3 0
1 241 0 4 0
1 246 0 6 0
1 253 0 2 0
1 256 0 2 0
1 259 0 2 0
1 262 0 1 0
1 263 0 2 0
1 266 0 2 0
1 269 0 2 0
1 272 0 2 0
1 275 0 2 0
1 278 0 2 0
1 281 0 2 0
1 284 0 2 0
1 287 0 2 0
1 290 0 3 0
1 294 0 2 0
1 297 0 3 0
1 301 0 3 0
1 305 0 3 0
1 309 0 3 0
1 313 0 2 0
1 316 0 2 0
1 319 0 2 0
1 322 0 2 0
1 325 0 2 0
1 328 0 2 0
1 331 0 2 0
1 334 0 2 0
1 337 0 2 0
1 340 0 2 0
1 343 0 2 0
1 346 0 2 0
1 349 0 2 0
1 352 0 2 0
1 355 0 2 0
3 398 1 0 1 220
3 400 1 0 1 221
3 401 1 0 1 222
0 405 7 1 2 1 3
0 408 5 1 1 230
3 419 1 0 1 254
3 420 1 0 1 255
0 425 5 1 1 262
3 456 1 0 1 291
3 457 1 0 1 292
3 458 1 0 1 293
0 485 7 1 4 310 306 302 298
0 486 5 1 1 405
3 487 5 0 1 45
3 488 5 0 1 133
3 489 5 0 1 83
3 490 5 0 1 97
3 491 5 0 1 70
3 492 5 0 1 121
3 493 5 0 1 58
3 494 5 0 1 109
0 495 7 1 3 2 15 238
0 496 1 2 1 239
0 499 7 1 2 38 38
0 500 1 2 1 223
0 503 1 2 1 9
0 506 1 2 1 10
0 509 1 11 1 228
0 521 1 11 1 235
0 533 5 3 1 242
0 537 5 5 1 247
0 543 7 1 2 12 248
0 544 7 2 4 134 84 98 46
0 547 7 2 4 122 59 110 71
0 550 1 11 1 229
0 562 1 11 1 236
0 574 5 3 1 257
0 578 5 3 1 260
0 582 1 11 1 320
0 594 1 11 1 323
0 606 5 1 1 329
0 607 5 1 1 332
0 608 5 1 1 335
0 609 5 1 1 338
0 610 5 1 1 341
0 611 5 1 1 344
0 612 5 1 1 353
0 613 1 11 1 321
0 625 1 11 1 324
0 637 1 5 1 17
0 643 1 6 1 18
0 650 5 1 1 356
0 651 7 3 2 7 240
0 655 5 3 1 264
0 659 5 3 1 267
0 663 5 3 1 270
0 667 5 3 1 273
0 671 5 3 1 276
0 675 5 3 1 279
0 679 5 3 1 282
0 683 5 3 1 285
0 687 5 5 1 288
0 693 1 5 1 30
0 699 1 5 1 31
0 705 5 5 1 295
0 711 5 3 1 299
0 715 5 3 1 303
0 719 5 3 1 307
0 723 5 3 1 311
0 727 5 2 1 314
0 730 5 2 1 317
0 733 5 1 1 347
0 734 5 1 1 350
0 735 1 2 1 261
0 738 1 2 1 258
0 741 1 2 1 265
0 744 1 2 1 271
0 747 1 2 1 268
0 750 1 2 1 277
0 753 1 2 1 274
0 756 1 2 1 283
0 759 1 2 1 280
0 762 1 2 1 289
0 765 1 2 1 286
0 768 1 2 1 296
0 771 1 2 1 304
0 774 1 2 1 300
0 777 1 2 1 312
0 780 1 2 1 308
0 783 1 2 1 318
0 786 1 2 1 315
3 792 5 0 1 485
3 799 5 0 1 495
0 800 5 2 1 499
3 805 1 0 1 360
0 900 6 1 2 333 606
0 901 6 1 2 330 607
0 902 6 1 2 339 608
0 903 6 1 2 336 609
0 904 6 1 2 345 610
0 905 6 1 2 342 611
0 998 6 1 2 351 733
0 999 6 1 2 348 734
3 1026 7 0 2 94 361
0 1027 7 1 2 326 511
3 1028 5 0 1 512
3 1029 6 0 2 232 513
0 1032 5 1 1 396
0 1033 5 1 1 399
0 1034 7 2 2 402 397
0 1037 1 4 1 362
0 1042 5 10 1 366
0 1053 5 10 1 377
0 1064 7 1 3 80 367 378
0 1065 7 1 3 68 368 379
0 1066 7 1 3 79 369 380
0 1067 7 1 3 78 370 381
0 1068 7 1 3 77 371 382
0 1069 7 1 2 13 391
0 1070 1 4 1 363
0 1075 5 10 1 403
0 1086 5 10 1 416
0 1097 7 1 3 76 404 417
0 1098 7 1 3 75 406 418
0 1099 7 1 3 74 407 421
0 1100 7 1 3 73 409 422
0 1101 7 1 3 72 410 423
0 1102 5 10 1 436
0 1113 5 10 1 447
0 1124 7 1 3 114 437 448
0 1125 7 1 3 113 438 449
0 1126 7 1 3 112 439 450
0 1127 7 1 3 111 440 451
0 1128 7 1 2 441 452
0 1129 6 3 2 900 901
0 1133 6 3 2 902 903
0 1137 6 2 2 904 905
0 1140 5 1 1 589
0 1141 6 1 2 590 612
0 1142 5 1 1 591
0 1143 5 1 1 593
0 1144 5 1 1 596
0 1145 5 1 1 598
0 1146 5 10 1 461
0 1157 5 10 1 472
0 1168 7 1 3 118 462 473
0 1169 7 1 3 107 463 474
0 1170 7 1 3 117 464 475
0 1171 7 1 3 116 465 476
0 1172 7 1 3 115 466 477
0 1173 5 4 1 483
0 1178 5 5 1 502
0 1184 5 1 1 616
0 1185 6 1 2 617 650
0 1186 5 1 1 618
0 1187 5 1 1 620
0 1188 5 1 1 622
0 1189 5 1 1 624
0 1190 1 4 1 364
0 1195 1 4 1 365
0 1200 5 4 1 549
0 1205 5 4 1 555
0 1210 5 1 1 585
0 1211 5 1 1 587
0 1212 5 1 1 600
0 1213 5 1 1 602
0 1214 5 1 1 604
0 1215 5 1 1 614
0 1216 6 2 2 998 999
0 1219 1 2 1 430
0 1222 1 2 1 433
0 1225 1 2 1 514
0 1228 1 2 1 517
0 1231 1 2 1 520
0 1234 1 2 1 524
0 1237 1 2 1 527
0 1240 1 2 1 530
0 1243 1 2 1 534
0 1246 1 2 1 538
0 1249 5 1 1 627
0 1250 5 1 1 629
0 1251 1 2 1 541
0 1254 1 2 1 560
0 1257 1 2 1 566
0 1260 1 2 1 569
0 1263 1 2 1 572
0 1266 1 2 1 576
3 1269 5 0 1 1027
0 1275 7 1 2 327 1032
0 1276 7 1 2 233 1033
3 1277 1 0 1 633
0 1302 3 1 2 1069 543
0 1351 6 1 2 354 1140
0 1352 6 1 2 595 1142
0 1353 6 1 2 592 1143
0 1354 6 1 2 599 1144
0 1355 6 1 2 597 1145
0 1395 6 1 2 357 1184
0 1396 6 1 2 621 1186
0 1397 6 1 2 619 1187
0 1398 6 1 2 626 1188
0 1399 6 1 2 623 1189
0 1422 6 1 2 588 1210
0 1423 6 1 2 586 1211
0 1424 6 1 2 603 1212
0 1425 6 1 2 601 1213
0 1426 6 1 2 615 1214
0 1427 6 1 2 605 1215
0 1440 6 1 2 630 1249
0 1441 6 1 2 628 1250
3 1448 5 0 1 634
0 1449 5 1 1 1275
0 1450 5 1 1 1276
0 1451 7 1 3 93 640 653
0 1452 7 1 3 55 372 654
0 1453 7 1 3 67 641 383
0 1454 7 1 3 81 642 656
0 1455 7 1 3 43 373 657
0 1456 7 1 3 56 644 384
0 1457 7 1 3 92 645 658
0 1458 7 1 3 54 374 660
0 1459 7 1 3 66 646 385
0 1460 7 1 3 91 647 661
0 1461 7 1 3 53 375 662
0 1462 7 1 3 65 648 386
0 1463 7 1 3 90 649 664
0 1464 7 1 3 52 376 665
0 1465 7 1 3 64 652 387
0 1466 7 1 3 89 672 685
0 1467 7 1 3 51 411 686
0 1468 7 1 3 63 673 424
0 1469 7 1 3 88 674 688
0 1470 7 1 3 50 412 689
0 1471 7 1 3 62 676 426
0 1472 7 1 3 87 677 690
0 1473 7 1 3 49 413 691
0 1474 7 1 2 678 427
0 1475 7 1 3 86 680 692
0 1476 7 1 3 48 414 694
0 1477 7 1 3 61 681 428
0 1478 7 1 3 85 682 695
0 1479 7 1 3 47 415 696
0 1480 7 1 3 60 684 429
0 1481 7 1 3 138 697 709
0 1482 7 1 3 102 442 710
0 1483 7 1 3 126 698 453
0 1484 7 1 3 137 700 712
0 1485 7 1 3 101 443 713
0 1486 7 1 3 125 701 454
0 1487 7 1 3 136 702 714
0 1488 7 1 3 100 444 716
0 1489 7 1 3 124 703 455
0 1490 7 1 3 135 704 717
0 1491 7 1 3 99 445 718
0 1492 7 1 3 123 706 459
0 1493 7 1 2 707 720
0 1494 7 1 2 446 721
0 1495 7 1 2 708 460
0 1496 5 2 1 722
0 1499 5 2 1 726
0 1502 6 3 2 1351 1141
0 1506 6 3 2 1352 1353
0 1510 6 2 2 1354 1355
0 1513 1 2 1 731
0 1516 1 2 1 732
0 1519 5 1 1 803
0 1520 5 1 1 806
0 1521 5 1 1 808
0 1522 5 1 1 810
0 1523 5 1 1 812
0 1524 5 1 1 814
0 1525 5 1 1 816
0 1526 5 1 1 818
0 1527 5 1 1 820
0 1528 5 1 1 822
0 1529 7 1 3 142 736 751
0 1530 7 1 3 106 467 752
0 1531 7 1 3 130 737 478
0 1532 7 1 3 131 739 754
0 1533 7 1 3 95 468 755
0 1534 7 1 3 119 740 479
0 1535 7 1 3 141 742 757
0 1536 7 1 3 105 469 758
0 1537 7 1 3 129 743 480
0 1538 7 1 3 140 745 760
0 1539 7 1 3 104 470 761
0 1540 7 1 3 128 746 481
0 1541 7 1 3 139 748 763
0 1542 7 1 3 103 471 764
0 1543 7 1 3 127 749 482
0 1544 7 1 2 19 766
0 1545 7 1 2 4 767
0 1546 7 1 2 20 769
0 1547 7 1 2 5 770
0 1548 7 1 2 21 772
0 1549 7 1 2 22 773
0 1550 7 1 2 23 775
0 1551 7 1 2 6 776
0 1552 7 1 2 24 778
0 1553 6 3 2 1395 1185
0 1557 6 3 2 1396 1397
0 1561 6 2 2 1398 1399
0 1564 7 1 2 25 790
0 1565 7 1 2 32 791
0 1566 7 1 2 26 793
0 1567 7 1 2 33 794
0 1568 7 1 2 27 795
0 1569 7 1 2 34 796
0 1570 7 1 2 35 797
0 1571 7 1 2 28 798
0 1572 5 1 1 824
0 1573 5 1 1 826
0 1574 5 1 1 828
0 1575 5 1 1 830
0 1576 5 1 1 832
0 1577 5 1 1 834
0 1578 6 2 2 1422 1423
0 1581 5 1 1 801
0 1582 6 2 2 1426 1427
0 1585 6 2 2 1424 1425
0 1588 6 2 2 1440 1441
0 1591 7 4 2 1449 1450
0 1596 3 3 4 1451 1452 1453 1064
0 1600 3 5 4 1454 1455 1456 1065
0 1606 3 5 4 1457 1458 1459 1066
0 1612 3 2 4 1460 1461 1462 1067
0 1615 3 3 4 1463 1464 1465 1068
0 1619 3 4 4 1466 1467 1468 1097
0 1624 3 3 4 1469 1470 1471 1098
0 1628 3 2 4 1472 1473 1474 1099
0 1631 3 2 4 1475 1476 1477 1100
0 1634 3 2 4 1478 1479 1480 1101
0 1637 3 4 4 1481 1482 1483 1124
0 1642 3 4 4 1484 1485 1486 1125
0 1647 3 3 4 1487 1488 1489 1126
0 1651 3 4 4 1490 1491 1492 1127
0 1656 3 3 4 1493 1494 1495 1128
0 1676 3 4 4 1532 1533 1534 1169
0 1681 3 4 4 1535 1536 1537 1170
0 1686 3 3 4 1538 1539 1540 1171
0 1690 3 2 4 1541 1542 1543 1172
0 1708 3 2 4 1529 1530 1531 1168
3 1726 1 0 1 868
0 1770 5 2 1 840
0 1773 5 2 1 843
0 1776 5 1 1 848
0 1777 5 1 1 850
0 1778 1 2 1 846
0 1781 1 2 1 847
0 1784 7 1 3 728 724 849
0 1785 7 1 3 838 836 851
0 1795 5 2 1 852
0 1798 5 2 1 855
0 1801 1 2 1 858
0 1804 1 2 1 859
0 1807 5 1 1 866
0 1808 5 1 1 860
0 1809 6 1 2 861 1581
0 1810 5 1 1 862
0 1811 5 1 1 864
0 1813 7 1 2 872 243
0 1814 7 1 2 880 244
0 1815 7 1 2 875 245
3 1816 5 0 1 913
3 1817 5 0 1 917
3 1818 5 0 1 909
3 1819 5 0 1 894
3 1820 5 0 1 890
3 1821 5 0 1 887
0 1822 7 1 4 358 225 36 869
0 1823 7 1 4 359 226 870 486
0 1824 1 2 1 873
0 1827 5 2 1 881
0 1830 7 1 2 876 392
0 1831 7 1 2 882 393
0 1832 7 1 2 891 249
0 1833 5 2 1 874
0 1836 5 4 1 877
0 1841 5 6 1 883
0 1848 1 3 1 885
0 1852 1 3 1 888
0 1856 1 6 1 892
0 1863 1 6 1 895
0 1870 1 4 1 897
0 1875 1 4 1 899
0 1880 1 4 1 907
0 1885 6 2 2 580 920
0 1888 6 2 2 583 924
0 1891 1 2 1 935
0 1894 7 2 2 910 425
0 1897 5 2 1 914
0 1908 7 1 3 837 729 1776
0 1909 7 1 3 725 839 1777
0 1910 7 1 2 878 484
0 1911 7 1 2 884 497
0 1912 7 1 2 886 498
0 1913 7 1 2 889 501
0 1914 7 1 2 893 504
0 1915 7 1 2 896 505
0 1916 7 1 2 898 507
0 1917 7 1 2 906 508
0 1918 7 1 2 908 510
0 1919 5 1 1 940
0 1928 7 1 2 927 551
0 1929 7 1 2 931 552
0 1930 7 1 2 936 553
0 1931 7 1 2 938 554
0 1932 7 1 2 911 556
0 1933 7 1 2 915 557
0 1934 7 1 2 918 558
0 1935 7 1 2 921 559
0 1936 1 2 1 879
0 1939 6 1 2 802 1808
0 1940 6 1 2 865 1810
0 1941 6 1 2 863 1811
0 1942 1 2 1 928
0 1945 1 2 1 937
0 1948 1 2 1 932
0 1951 1 2 1 912
0 1954 1 2 1 939
0 1957 1 2 1 919
0 1960 1 2 1 916
0 1963 1 2 1 925
0 1966 1 2 1 922
3 1969 3 0 2 388 1815
3 1970 5 0 1 1822
3 1971 5 0 1 1823
3 2010 1 0 1 974
3 2012 1 0 1 977
3 2014 1 0 1 980
3 2016 1 0 1 986
3 2018 1 0 1 992
3 2020 1 0 1 996
3 2022 1 0 1 1002
0 2028 5 1 1 946
0 2029 5 1 1 948
0 2030 4 1 2 1908 1784
0 2031 4 1 2 1909 1785
0 2032 7 1 3 844 841 947
0 2033 7 1 3 944 942 949
0 2034 3 1 2 1571 1935
0 2040 5 1 1 954
0 2041 5 1 1 956
0 2042 7 1 3 856 853 955
0 2043 7 1 3 952 950 957
0 2046 6 2 2 1939 1809
0 2049 6 2 2 1940 1941
0 2052 3 2 2 1544 1910
0 2055 3 2 2 1545 1911
0 2058 3 2 2 1546 1912
0 2061 3 2 2 1547 1913
0 2064 3 2 2 1548 1914
0 2067 3 2 2 1549 1915
0 2070 3 2 2 1550 1916
0 2073 3 2 2 1551 1917
0 2076 3 2 2 1552 1918
0 2079 3 2 2 1564 1928
0 2095 3 2 2 1565 1929
0 2098 3 2 2 1566 1930
0 2101 3 2 2 1567 1931
0 2104 3 2 2 1568 1932
0 2107 3 2 2 1569 1933
0 2110 3 2 2 1570 1934
0 2113 7 5 3 1014 1012 41
0 2119 5 1 1 1013
0 2120 6 4 2 408 960
0 2125 7 1 2 958 394
0 2126 7 1 2 978 250
0 2127 7 1 2 975 395
0 2128 5 6 1 976
0 2135 5 5 1 979
0 2141 5 2 1 987
0 2144 5 2 1 993
0 2147 5 2 1 997
0 2150 5 2 1 1003
0 2153 7 1 2 581 1006
0 2154 7 1 2 1007 923
0 2155 7 1 2 584 1008
0 2156 7 1 2 1009 926
0 2157 7 1 3 943 845 2028
0 2158 7 1 3 842 945 2029
0 2171 5 1 1 1018
0 2172 6 1 2 1019 1919
0 2173 5 1 1 1020
0 2174 5 1 1 1022
0 2175 5 1 1 1024
0 2176 5 1 1 1030
0 2177 7 1 3 951 857 2040
0 2178 7 1 3 854 953 2041
0 2185 1 2 1 964
0 2188 1 2 1 962
0 2191 1 2 1 968
0 2194 5 2 1 981
0 2197 5 2 1 961
0 2200 5 1 1 1016
0 2201 1 2 1 965
0 2204 1 2 1 963
0 2207 1 2 1 969
0 2210 1 2 1 959
0 2213 1 2 1 970
0 2216 1 2 1 971
0 2219 6 2 2 2031 2030
0 2234 5 1 1 1035
0 2235 5 1 1 1038
0 2236 5 1 1 1040
0 2237 5 1 1 1043
0 2250 7 2 3 42 1015 2119
0 2266 3 2 2 1831 2126
0 2269 3 2 2 2127 1832
0 2291 3 2 2 2153 2154
0 2294 3 2 2 2155 2156
0 2297 4 1 2 2157 2032
0 2298 4 1 2 2158 2033
0 2300 5 1 1 1045
0 2301 5 1 1 1047
0 2302 6 1 2 1049 1519
0 2303 5 1 1 1050
0 2304 6 1 2 1051 1520
0 2305 5 1 1 1052
0 2306 6 1 2 1054 1521
0 2307 5 1 1 1055
0 2308 6 1 2 1056 1522
0 2309 5 1 1 1057
0 2310 6 1 2 1058 1523
0 2311 5 1 1 1059
0 2312 6 1 2 1060 1524
0 2313 5 1 1 1061
0 2314 6 1 2 1062 1525
0 2315 5 1 1 1063
0 2316 6 1 2 1071 1526
0 2317 5 1 1 1072
0 2318 6 1 2 1073 1527
0 2319 5 1 1 1074
0 2320 6 1 2 1076 1528
0 2321 5 1 1 1077
0 2322 6 1 2 941 2171
0 2323 6 1 2 1023 2173
0 2324 6 1 2 1021 2174
0 2325 6 1 2 1031 2175
0 2326 6 1 2 1025 2176
0 2327 4 1 2 2177 2042
0 2328 4 1 2 2178 2043
0 2329 6 1 2 1078 1572
0 2330 5 1 1 1079
0 2331 6 1 2 1080 1573
0 2332 5 1 1 1081
0 2333 6 1 2 1082 1574
0 2334 5 1 1 1083
0 2335 6 1 2 1084 1575
0 2336 5 1 1 1085
0 2337 6 1 2 1087 1576
0 2338 5 1 1 1088
0 2339 6 1 2 1089 1577
0 2340 5 1 1 1090
0 2354 6 1 2 1039 2234
0 2355 6 1 2 1036 2235
0 2356 6 1 2 1044 2236
0 2357 6 1 2 1041 2237
0 2358 7 1 2 1096 389
0 2359 5 2 1 1091
0 2364 5 1 1 1132
0 2365 5 1 1 1135
0 2366 5 1 1 1138
0 2367 5 1 1 1147
0 2368 1 3 1 1103
0 2372 5 1 1 1151
0 2373 5 1 1 1153
0 2374 5 1 1 1155
0 2375 5 1 1 1158
0 2376 5 1 1 1160
0 2377 5 4 1 1092
0 2382 1 3 1 1093
0 2386 7 1 2 1104 251
3 2387 1 0 1 1174
3 2388 1 0 1 1175
3 2389 1 0 1 1176
3 2390 1 0 1 1177
0 2391 1 3 1 1094
0 2395 5 4 1 1095
0 2400 6 1 2 1164 2300
0 2403 5 1 1 1162
0 2406 5 1 1 1165
0 2407 6 1 2 804 2303
0 2408 6 1 2 807 2305
0 2409 6 1 2 809 2307
0 2410 6 1 2 811 2309
0 2411 6 1 2 813 2311
0 2412 6 1 2 815 2313
0 2413 6 1 2 817 2315
0 2414 6 1 2 819 2317
0 2415 6 1 2 821 2319
0 2416 6 1 2 823 2321
0 2417 6 3 2 2322 2172
0 2421 6 3 2 2323 2324
0 2425 6 2 2 2325 2326
0 2428 6 1 2 825 2330
0 2429 6 1 2 827 2332
0 2430 6 1 2 829 2334
0 2431 6 1 2 831 2336
0 2432 6 1 2 833 2338
0 2433 6 1 2 835 2340
0 2434 1 2 1 1106
0 2437 1 2 1 1112
0 2440 1 2 1 1120
0 2443 1 2 1 1118
0 2446 1 2 1 1130
0 2449 1 2 1 1122
0 2452 5 1 1 1149
0 2453 6 1 2 1150 2200
0 2454 1 2 1 1107
0 2457 1 2 1 1121
0 2460 1 2 1 1119
0 2463 1 2 1 1131
0 2466 1 2 1 1123
0 2469 5 2 1 1105
0 2472 1 2 1 1108
0 2475 1 2 1 1114
0 2478 1 2 1 1109
0 2481 1 2 1 1115
0 2484 6 2 2 2298 2297
0 2487 6 2 2 2356 2357
0 2490 6 2 2 2354 2355
0 2493 6 2 2 2328 2327
3 2496 3 0 2 2358 1814
0 2503 6 1 2 1136 2364
0 2504 6 1 2 1134 2365
0 2510 6 1 2 1154 2372
0 2511 6 1 2 1152 2373
0 2521 3 2 2 1830 2386
0 2528 6 1 2 1046 2406
0 2531 5 2 1 1179
0 2534 5 2 1 1181
0 2537 1 2 1 1166
0 2540 1 2 1 1167
0 2544 6 1 2 2302 2407
0 2545 6 1 2 2304 2408
0 2546 6 1 2 2306 2409
0 2547 6 1 2 2308 2410
0 2548 6 1 2 2310 2411
0 2549 6 1 2 2312 2412
0 2550 6 1 2 2314 2413
0 2551 6 1 2 2316 2414
0 2552 6 1 2 2318 2415
0 2553 6 1 2 2320 2416
0 2563 6 1 2 2329 2428
0 2564 6 1 2 2331 2429
0 2565 6 1 2 2333 2430
0 2566 6 1 2 2335 2431
0 2567 6 1 2 2337 2432
0 2568 6 1 2 2339 2433
0 2579 6 1 2 1017 2452
0 2603 1 3 1 1183
0 2607 7 1 2 1004 1196
0 2608 7 1 2 929 1197
0 2609 7 1 2 933 1198
0 2610 7 1 2 1010 1199
0 2611 7 1 2 982 1201
0 2612 7 1 2 988 1202
0 2613 6 3 2 2503 2504
0 2617 5 1 1 1232
0 2618 6 1 2 1233 2366
0 2619 6 1 2 1235 2367
0 2620 5 1 1 1236
0 2621 5 2 1 1192
0 2624 6 3 2 2510 2511
0 2628 5 1 1 1252
0 2629 6 1 2 1253 2374
0 2630 5 1 1 1270
0 2631 7 1 2 983 1204
0 2632 7 1 2 989 1206
0 2633 7 1 2 1005 1208
0 2634 7 1 2 930 1209
0 2635 7 1 2 934 1217
0 2636 7 1 2 1011 1218
0 2638 5 4 1 1203
3 2643 1 0 1 1289
3 2644 1 0 1 1290
0 2645 5 1 1 1272
0 2646 5 4 1 1207
0 2652 6 1 2 2528 2400
0 2655 5 1 1 1274
0 2656 5 1 1 1279
0 2659 1 3 1 1191
0 2663 5 1 1 1281
0 2664 6 1 2 1282 2301
0 2665 5 1 1 2553
0 2666 5 1 1 2552
0 2667 5 1 1 2551
0 2668 5 1 1 2550
0 2669 5 1 1 2549
0 2670 5 1 1 2548
0 2671 5 1 1 2547
0 2672 5 1 1 2546
0 2673 5 1 1 2545
0 2674 5 1 1 2544
0 2675 5 1 1 2568
0 2676 5 1 1 2567
0 2677 5 1 1 2566
0 2678 5 1 1 2565
0 2679 5 1 1 2564
0 2680 5 1 1 2563
0 2681 5 2 1 1220
0 2684 5 2 1 1224
0 2687 1 2 1 1229
0 2690 1 2 1 1230
0 2693 5 1 1 1287
0 2694 6 1 2 1288 1807
0 2695 5 1 1 1238
0 2696 5 1 1 1241
0 2697 5 1 1 1244
0 2698 5 1 1 1247
0 2699 5 1 1 1255
0 2700 5 1 1 1258
0 2701 5 1 1 1261
0 2702 5 1 1 1264
0 2703 6 2 2 2579 2453
0 2706 5 1 1 1267
0 2707 5 1 1 1283
0 2708 5 1 1 1285
0 2709 7 1 2 1182 1293
0 2710 7 1 2 1180 1291
0 2719 6 1 2 1139 2617
0 2720 6 1 2 1148 2620
0 2726 6 1 2 1156 2628
0 2729 1 4 1 1295
0 2738 1 4 1 1296
0 2743 5 1 1 2652
0 2747 6 1 2 1048 2663
0 2748 7 1 5 2665 2666 2667 2668 2669
0 2749 7 1 5 2670 2671 2672 2673 2674
0 2750 7 1 2 2034 2675
0 2751 7 1 5 2676 2677 2678 2679 2680
0 2760 6 1 2 867 2693
0 2761 1 4 1 1297
0 2766 1 4 1 1298
0 2771 6 1 2 1242 2695
0 2772 6 1 2 1239 2696
0 2773 6 1 2 1248 2697
0 2774 6 1 2 1245 2698
0 2775 6 1 2 1259 2699
0 2776 6 1 2 1256 2700
0 2777 6 1 2 1265 2701
0 2778 6 1 2 1262 2702
0 2781 6 1 2 1286 2707
0 2782 6 1 2 1284 2708
0 2783 3 1 2 2709 1294
0 2784 3 1 2 2710 1292
0 2789 7 1 2 984 1311
0 2790 7 1 2 990 1312
0 2791 7 1 2 994 1313
0 2792 7 1 2 1000 1314
0 2793 5 2 1 1303
0 2796 6 3 2 2719 2618
0 2800 6 2 2 2619 2720
0 2803 5 2 1 1308
0 2806 6 2 2 2726 2629
0 2809 7 1 2 985 1315
0 2810 7 1 2 991 1316
0 2811 7 1 2 995 1317
0 2812 7 1 2 1001 1318
0 2817 7 2 2 2743 14
0 2820 1 5 1 1299
0 2826 6 2 2 2747 2664
0 2829 7 1 2 2748 2749
0 2830 7 1 2 2750 2751
0 2831 1 5 1 1319
0 2837 5 1 1 1326
0 2838 5 1 1 1328
0 2839 7 1 3 1226 1221 1327
0 2840 7 1 3 1324 1322 1329
0 2841 6 2 2 2760 2694
0 2844 1 5 1 1300
0 2854 1 4 1 1301
0 2859 1 5 1 1320
0 2869 1 4 1 1321
0 2874 6 2 2 2773 2774
0 2877 6 2 2 2771 2772
0 2880 5 1 1 1330
0 2881 6 1 2 1331 2706
0 2882 6 2 2 2777 2778
0 2885 6 2 2 2775 2776
0 2888 6 2 2 2781 2782
3 2891 6 0 2 2783 2784
0 2894 7 1 2 2607 1332
0 2895 7 1 2 2608 1333
0 2896 7 1 2 2609 1334
0 2897 7 1 2 2610 1335
0 2898 3 1 2 2789 2611
0 2899 3 1 2 2790 2612
0 2900 7 1 2 2791 635
0 2901 7 1 2 2792 636
0 2914 3 1 2 2809 2631
0 2915 3 1 2 2810 2632
0 2916 7 1 2 2811 666
0 2917 7 1 2 2812 668
0 2918 7 1 2 2633 1336
0 2919 7 1 2 2634 1337
0 2920 7 1 2 2635 1338
0 2921 7 1 2 2636 1339
3 2925 1 0 1 1364
0 2931 7 2 3 2829 2830 1302
0 2938 7 1 3 1323 1227 2837
0 2939 7 1 3 1223 1325 2838
0 2963 6 1 2 1268 2880
3 2970 5 0 1 1378
3 2971 5 0 1 1371
0 2972 5 2 1 2894
0 2975 5 2 1 2895
0 2978 5 2 1 2896
0 2981 5 2 1 2897
0 2984 7 1 2 2898 638
0 2985 7 1 2 2899 639
0 2986 5 2 1 2900
0 2989 5 2 1 2901
0 2992 5 2 1 1350
0 2995 1 2 1 1358
0 2998 1 2 1 1359
0 3001 1 2 1 1362
0 3004 1 2 1 1363
0 3007 7 1 2 431 1366
0 3008 7 1 2 2914 669
0 3009 7 1 2 2915 670
0 3010 5 2 1 2916
0 3013 5 2 1 2917
0 3016 5 2 1 2918
0 3019 5 2 1 2919
0 3022 5 2 1 2920
0 3025 5 2 1 2921
0 3028 5 1 1 1365
0 3029 7 1 2 432 1373
0 3030 5 4 1 1367
0 3035 7 1 2 434 1368
0 3036 7 1 2 515 1369
0 3037 7 1 2 518 1370
3 3038 1 0 1 1413
0 3039 5 4 1 1374
0 3044 7 1 2 435 1375
0 3045 7 1 2 516 1376
0 3046 7 1 2 519 1377
0 3047 4 1 2 2938 2839
0 3048 4 1 2 2939 2840
0 3049 5 1 1 1411
0 3050 5 2 1 1380
0 3053 7 1 2 522 1381
0 3054 7 1 2 525 1382
0 3055 7 1 2 528 1383
0 3056 7 1 2 531 1384
0 3057 7 1 2 535 1385
0 3058 7 1 2 539 1386
0 3059 7 1 2 542 1387
0 3060 7 1 2 561 1388
0 3061 5 2 1 1389
0 3064 7 1 2 523 1390
0 3065 7 1 2 526 1391
0 3066 7 1 2 529 1392
0 3067 7 1 2 532 1393
0 3068 7 1 2 536 1394
0 3069 7 1 2 540 1400
0 3070 7 1 2 545 1401
0 3071 7 1 2 563 1402
0 3072 5 1 1 1403
0 3073 5 1 1 1405
0 3074 5 1 1 1407
0 3075 5 1 1 1409
0 3076 6 2 2 2881 2963
3 3079 5 0 1 1414
0 3088 5 2 1 2984
0 3091 5 2 1 2985
0 3110 5 2 1 3008
0 3113 5 2 1 3009
0 3137 7 2 2 3055 779
0 3140 7 2 2 3056 781
0 3143 7 2 2 3057 1340
0 3146 7 2 2 3058 1341
0 3149 7 2 2 3059 1342
0 3152 7 2 2 3060 1343
0 3157 7 2 2 3066 785
0 3160 7 2 2 3067 787
0 3163 7 2 2 3068 1344
0 3166 7 2 2 3069 1345
0 3169 7 2 2 3070 1346
0 3172 7 2 2 3071 1347
0 3175 6 1 2 1406 3072
0 3176 6 1 2 1404 3073
0 3177 6 1 2 1410 3074
0 3178 6 1 2 1408 3075
0 3180 6 2 2 3048 3047
0 3187 5 1 1 1435
0 3188 5 1 1 1437
0 3189 5 1 1 1439
0 3190 5 1 1 1443
0 3191 7 1 3 1356 1304 1436
0 3192 7 1 3 1433 1348 1438
0 3193 7 1 3 1309 1193 1442
0 3194 7 1 3 1360 1306 1444
0 3195 6 1 2 1560 2375
0 3196 5 1 1 1562
0 3197 7 1 2 546 1509
0 3208 7 1 2 548 1515
0 3215 7 1 2 564 1511
0 3216 7 1 2 567 1512
0 3217 7 1 2 570 1514
0 3218 7 1 2 565 1517
0 3219 7 1 2 568 1518
0 3220 7 1 2 571 1554
0 3222 7 1 2 573 1555
0 3223 7 1 2 577 1556
0 3230 7 1 2 575 1558
0 3231 7 1 2 579 1559
0 3238 6 2 2 3175 3176
0 3241 6 2 2 3177 3178
0 3244 1 2 1 1421
0 3247 1 2 1 1419
0 3250 1 2 1 1417
0 3253 1 2 1 1415
0 3256 1 2 1 1431
0 3259 1 2 1 1429
0 3262 1 2 1 1507
0 3265 1 2 1 1504
0 3268 1 2 1 1501
0 3271 1 2 1 1498
0 3274 1 2 1 1447
0 3277 1 2 1 1445
0 3281 7 1 3 1349 1357 3187
0 3282 7 1 3 1305 1434 3188
0 3283 7 1 3 1307 1310 3189
0 3284 7 1 3 1194 1361 3190
0 3286 6 1 2 1159 3196
0 3288 3 1 2 3197 3007
0 3289 6 1 2 1621 3049
0 3291 7 1 2 1603 1428
0 3293 7 1 2 1601 1420
0 3295 7 1 2 1598 1418
0 3296 7 1 2 1416 1595
0 3299 7 1 2 1593 1432
0 3301 7 1 2 1590 1430
0 3302 3 1 2 3208 3029
0 3304 7 1 2 1618 1508
0 3306 7 1 2 1616 1505
0 3308 7 1 2 1613 1503
0 3309 7 1 2 1500 1610
0 3312 7 1 2 1608 1497
0 3314 7 1 2 1605 1446
0 3315 3 2 2 3215 3035
0 3318 3 2 2 3216 3036
0 3321 3 2 2 3217 3037
0 3324 3 2 2 3218 3044
0 3327 3 2 2 3219 3045
0 3330 3 2 2 3220 3046
0 3333 5 1 1 1622
0 3334 3 1 2 3222 3053
0 3335 3 1 2 3223 3054
0 3336 3 1 2 3230 3064
0 3337 3 1 2 3231 3065
0 3340 1 2 1 1604
0 3344 1 2 1 1602
0 3348 1 2 1 1599
0 3352 1 2 1 1597
0 3356 1 2 1 1594
0 3360 1 2 1 1592
0 3364 1 2 1 1580
0 3367 1 2 1 1563
0 3370 1 2 1 1620
0 3374 1 2 1 1617
0 3378 1 2 1 1614
0 3382 1 2 1 1611
0 3386 1 2 1 1609
0 3390 1 2 1 1607
0 3394 1 2 1 1587
0 3397 1 2 1 1584
0 3400 6 1 2 3195 3286
0 3401 4 1 2 3281 3191
0 3402 4 1 2 3282 3192
0 3403 4 1 2 3283 3193
0 3404 4 1 2 3284 3194
0 3405 5 1 1 1623
0 3406 5 1 1 1626
0 3409 7 1 2 3288 966
0 3410 6 1 2 1412 3333
0 3412 5 1 1 1629
0 3414 5 1 1 1632
0 3416 5 1 1 1635
0 3418 5 1 1 1638
0 3420 5 1 1 1640
0 3422 5 1 1 1643
0 3428 7 1 2 3302 967
0 3430 5 1 1 1645
0 3432 5 1 1 1648
0 3434 5 1 1 1650
0 3436 5 1 1 1653
0 3438 5 1 1 1655
0 3440 5 1 1 1658
0 3450 7 2 2 3334 782
0 3453 7 2 2 3335 784
0 3456 7 2 2 3336 788
0 3459 7 2 2 3337 789
0 3478 7 1 2 3400 390
0 3479 7 1 2 1662 1110
0 3480 7 1 2 1660 972
0 3481 6 1 2 3410 3289
0 3482 5 1 1 1672
0 3483 6 1 2 1673 3412
0 3484 5 1 1 1674
0 3485 6 1 2 1675 3414
0 3486 5 1 1 1677
0 3487 6 1 2 1678 3416
0 3488 5 1 1 1679
0 3489 6 1 2 1680 3418
0 3490 5 1 1 1682
0 3491 6 1 2 1683 3420
0 3492 5 1 1 1684
0 3493 6 1 2 1685 3422
0 3494 5 1 1 1687
0 3496 5 1 1 1689
0 3498 7 1 2 1664 1116
0 3499 7 1 2 1668 1111
0 3500 7 1 2 1666 973
0 3501 5 1 1 1692
0 3502 6 1 2 1693 3430
0 3503 5 1 1 1694
0 3504 6 1 2 1695 3432
0 3505 5 1 1 1696
0 3506 6 1 2 1697 3434
0 3507 5 1 1 1698
0 3508 6 1 2 1699 3436
0 3509 5 1 1 1700
0 3510 6 1 2 1701 3438
0 3511 5 1 1 1702
0 3512 6 1 2 1703 3440
0 3513 5 1 1 1704
0 3515 5 1 1 1706
0 3517 7 1 2 1670 1117
0 3522 6 2 2 3402 3401
0 3525 6 2 2 3404 3403
0 3528 1 2 1 1663
0 3531 1 2 1 1661
0 3534 1 2 1 1665
0 3537 1 2 1 1669
0 3540 1 2 1 1667
0 3543 1 2 1 1671
3 3546 3 0 2 3478 1813
0 3551 5 1 1 3481
0 3552 6 1 2 1630 3482
0 3553 6 1 2 1633 3484
0 3554 6 1 2 1636 3486
0 3555 6 1 2 1639 3488
0 3556 6 1 2 1641 3490
0 3557 6 1 2 1644 3492
0 3558 7 1 2 1711 1583
0 3559 7 1 2 1709 1579
0 3563 6 1 2 1646 3501
0 3564 6 1 2 1649 3503
0 3565 6 1 2 1652 3505
0 3566 6 1 2 1654 3507
0 3567 6 1 2 1657 3509
0 3568 6 1 2 1659 3511
0 3569 7 1 2 1715 1589
0 3570 7 1 2 1713 1586
0 3576 1 2 1 1712
0 3579 1 2 1 1710
0 3585 1 2 1 1716
0 3588 1 2 1 1714
0 3592 5 1 1 1717
0 3593 6 1 2 1718 3405
0 3594 5 1 1 1719
0 3595 6 1 2 1720 3406
0 3596 5 1 1 1721
0 3597 6 1 2 1722 2630
0 3598 6 1 2 1723 2376
0 3599 5 1 1 1724
0 3600 7 2 2 3551 631
0 3603 6 4 2 3552 3483
0 3608 6 3 2 3553 3485
0 3612 6 2 2 3554 3487
0 3615 6 1 2 3555 3489
0 3616 6 5 2 3556 3491
0 3622 6 4 2 3557 3493
0 3629 5 1 1 1725
0 3630 6 1 2 1727 2645
0 3631 5 1 1 1728
0 3632 6 1 2 1729 2655
0 3633 6 1 2 1730 2403
0 3634 5 1 1 1731
0 3635 6 4 2 3563 3502
0 3640 6 3 2 3564 3504
0 3644 6 2 2 3565 3506
0 3647 6 1 2 3566 3508
0 3648 6 5 2 3567 3510
0 3654 6 4 2 3568 3512
0 3661 5 1 1 1732
0 3662 6 1 2 1733 2656
0 3667 6 1 2 1625 3592
0 3668 6 1 2 1627 3594
0 3669 6 1 2 1271 3596
0 3670 6 1 2 1161 3599
3 3671 1 0 1 1742
0 3691 5 1 1 1734
0 3692 6 1 2 1735 3494
0 3693 5 1 1 1736
0 3694 6 1 2 1737 3496
0 3695 6 1 2 1273 3629
0 3696 6 1 2 1278 3631
0 3697 6 1 2 1163 3634
0 3716 5 1 1 1738
0 3717 6 1 2 1739 3513
0 3718 5 1 1 1740
0 3719 6 1 2 1741 3515
0 3720 6 1 2 1280 3661
0 3721 6 1 2 3667 3593
0 3722 6 1 2 3668 3595
0 3723 6 2 2 3669 3597
0 3726 6 1 2 3670 3598
0 3727 5 1 1 1743
0 3728 6 1 2 1688 3691
0 3729 6 1 2 1691 3693
0 3730 6 1 2 3695 3630
0 3731 7 1 4 1748 3615 1751 1744
0 3732 7 1 2 1745 3293
0 3733 7 1 3 1749 1746 3295
0 3734 7 1 4 1752 1747 3296 1750
0 3735 7 1 2 1753 3301
0 3736 7 1 3 1758 1754 3558
0 3737 6 2 2 3696 3632
0 3740 6 1 2 3697 3633
0 3741 6 1 2 1705 3716
0 3742 6 1 2 1707 3718
0 3743 6 1 2 3720 3662
0 3744 7 1 4 1766 3647 1769 1762
0 3745 7 1 2 1763 3306
0 3746 7 1 3 1767 1764 3308
0 3747 7 1 4 1771 1765 3309 1768
0 3748 7 1 2 1772 3314
0 3749 7 1 3 1782 1774 3569
0 3750 5 1 1 3721
0 3753 7 1 2 3722 252
0 3754 6 3 2 3728 3692
0 3758 6 2 2 3729 3694
0 3761 5 1 1 3731
0 3762 3 2 4 3291 3732 3733 3734
0 3767 6 3 2 3741 3717
0 3771 6 2 2 3742 3719
0 3774 5 1 1 3744
0 3775 3 2 4 3304 3745 3746 3747
0 3778 7 1 2 1788 3480
0 3779 7 1 3 3726 1789 3409
0 3780 3 2 2 2125 3753
0 3790 7 2 2 3750 632
0 3793 7 1 2 1790 3500
0 3794 7 1 3 3740 1791 3428
0 3802 3 1 3 3479 3778 3779
3 3803 1 0 1 1828
3 3804 1 0 1 1829
0 3805 5 1 1 1799
0 3806 7 1 5 1759 3730 1792 1755 1796
0 3807 7 1 4 1793 1756 3559 1760
0 3808 7 1 5 1797 1794 1757 3498 1761
3 3809 1 0 1 1834
0 3811 3 1 3 3499 3793 3794
0 3812 5 1 1 1825
0 3813 7 1 5 1783 3743 1802 1775 1806
0 3814 7 1 4 1803 1779 3570 1786
0 3815 7 1 5 1812 1805 1780 3517 1787
0 3816 3 1 5 3299 3735 3736 3807 3808
0 3817 7 1 2 3806 3802
0 3818 6 1 2 3805 3761
0 3819 5 1 1 1835
0 3820 3 1 5 3312 3748 3749 3814 3815
0 3821 7 1 2 3813 3811
0 3822 6 1 2 3812 3774
0 3823 3 2 2 3816 3817
0 3826 7 1 3 3727 3819 1379
0 3827 3 2 2 3820 3821
0 3834 5 1 1 1837
0 3835 7 1 2 3818 1838
0 3836 5 1 1 1839
0 3837 7 1 2 3822 1840
0 3838 7 1 2 1800 3834
0 3839 7 1 2 1826 3836
0 3840 3 2 2 3838 3835
0 3843 3 3 2 3839 3837
3 3851 1 0 1 1844
0 3852 6 2 2 1845 1842
0 3857 7 1 2 1846 1847
0 3858 7 1 2 1849 1843
0 3859 3 2 2 3857 3858
0 3864 5 2 1 1850
0 3869 7 1 2 1851 1853
0 3870 3 2 2 3869 1854
3 3875 5 0 1 1855
0 3876 7 1 3 1372 3028 1857
0 3877 7 2 3 3826 3876 871
3 3881 1 0 1 1858
3 3882 5 0 1 1859
2 9 1 8
2 10 1 8
2 12 1 11
2 13 1 11
2 17 1 16
2 18 1 16
2 30 1 29
2 31 1 29
2 38 1 37
2 39 1 37
2 41 1 40
2 42 1 40
2 45 1 44
2 46 1 44
2 58 1 57
2 59 1 57
2 70 1 69
2 71 1 69
2 83 1 82
2 84 1 82
2 97 1 96
2 98 1 96
2 109 1 108
2 110 1 108
2 121 1 120
2 122 1 120
2 133 1 132
2 134 1 132
2 220 1 219
2 221 1 219
2 222 1 219
2 223 1 219
2 225 1 224
2 226 1 224
2 228 1 227
2 229 1 227
2 232 1 231
2 233 1 231
2 235 1 234
2 236 1 234
2 238 1 237
2 239 1 237
2 240 1 237
2 242 1 241
2 243 1 241
2 244 1 241
2 245 1 241
2 247 1 246
2 248 1 246
2 249 1 246
2 250 1 246
2 251 1 246
2 252 1 246
2 254 1 253
2 255 1 253
2 257 1 256
2 258 1 256
2 260 1 259
2 261 1 259
2 264 1 263
2 265 1 263
2 267 1 266
2 268 1 266
2 270 1 269
2 271 1 269
2 273 1 272
2 274 1 272
2 276 1 275
2 277 1 275
2 279 1 278
2 280 1 278
2 282 1 281
2 283 1 281
2 285 1 284
2 286 1 284
2 288 1 287
2 289 1 287
2 291 1 290
2 292 1 290
2 293 1 290
2 295 1 294
2 296 1 294
2 298 1 297
2 299 1 297
2 300 1 297
2 302 1 301
2 303 1 301
2 304 1 301
2 306 1 305
2 307 1 305
2 308 1 305
2 310 1 309
2 311 1 309
2 312 1 309
2 314 1 313
2 315 1 313
2 317 1 316
2 318 1 316
2 320 1 319
2 321 1 319
2 323 1 322
2 324 1 322
2 326 1 325
2 327 1 325
2 329 1 328
2 330 1 328
2 332 1 331
2 333 1 331
2 335 1 334
2 336 1 334
2 338 1 337
2 339 1 337
2 341 1 340
2 342 1 340
2 344 1 343
2 345 1 343
2 347 1 346
2 348 1 346
2 350 1 349
2 351 1 349
2 353 1 352
2 354 1 352
2 356 1 355
2 357 1 355
2 358 1 496
2 359 1 496
2 360 1 500
2 361 1 500
2 362 1 503
2 363 1 503
2 364 1 506
2 365 1 506
2 366 1 509
2 367 1 509
2 368 1 509
2 369 1 509
2 370 1 509
2 371 1 509
2 372 1 509
2 373 1 509
2 374 1 509
2 375 1 509
2 376 1 509
2 377 1 521
2 378 1 521
2 379 1 521
2 380 1 521
2 381 1 521
2 382 1 521
2 383 1 521
2 384 1 521
2 385 1 521
2 386 1 521
2 387 1 521
2 388 1 533
2 389 1 533
2 390 1 533
2 391 1 537
2 392 1 537
2 393 1 537
2 394 1 537
2 395 1 537
2 396 1 544
2 397 1 544
2 399 1 547
2 402 1 547
2 403 1 550
2 404 1 550
2 406 1 550
2 407 1 550
2 409 1 550
2 410 1 550
2 411 1 550
2 412 1 550
2 413 1 550
2 414 1 550
2 415 1 550
2 416 1 562
2 417 1 562
2 418 1 562
2 421 1 562
2 422 1 562
2 423 1 562
2 424 1 562
2 426 1 562
2 427 1 562
2 428 1 562
2 429 1 562
2 430 1 574
2 431 1 574
2 432 1 574
2 433 1 578
2 434 1 578
2 435 1 578
2 436 1 582
2 437 1 582
2 438 1 582
2 439 1 582
2 440 1 582
2 441 1 582
2 442 1 582
2 443 1 582
2 444 1 582
2 445 1 582
2 446 1 582
2 447 1 594
2 448 1 594
2 449 1 594
2 450 1 594
2 451 1 594
2 452 1 594
2 453 1 594
2 454 1 594
2 455 1 594
2 459 1 594
2 460 1 594
2 461 1 613
2 462 1 613
2 463 1 613
2 464 1 613
2 465 1 613
2 466 1 613
2 467 1 613
2 468 1 613
2 469 1 613
2 470 1 613
2 471 1 613
2 472 1 625
2 473 1 625
2 474 1 625
2 475 1 625
2 476 1 625
2 477 1 625
2 478 1 625
2 479 1 625
2 480 1 625
2 481 1 625
2 482 1 625
2 483 1 637
2 484 1 637
2 497 1 637
2 498 1 637
2 501 1 637
2 502 1 643
2 504 1 643
2 505 1 643
2 507 1 643
2 508 1 643
2 510 1 643
2 511 1 651
2 512 1 651
2 513 1 651
2 514 1 655
2 515 1 655
2 516 1 655
2 517 1 659
2 518 1 659
2 519 1 659
2 520 1 663
2 522 1 663
2 523 1 663
2 524 1 667
2 525 1 667
2 526 1 667
2 527 1 671
2 528 1 671
2 529 1 671
2 530 1 675
2 531 1 675
2 532 1 675
2 534 1 679
2 535 1 679
2 536 1 679
2 538 1 683
2 539 1 683
2 540 1 683
2 541 1 687
2 542 1 687
2 545 1 687
2 546 1 687
2 548 1 687
2 549 1 693
2 551 1 693
2 552 1 693
2 553 1 693
2 554 1 693
2 555 1 699
2 556 1 699
2 557 1 699
2 558 1 699
2 559 1 699
2 560 1 705
2 561 1 705
2 563 1 705
2 564 1 705
2 565 1 705
2 566 1 711
2 567 1 711
2 568 1 711
2 569 1 715
2 570 1 715
2 571 1 715
2 572 1 719
2 573 1 719
2 575 1 719
2 576 1 723
2 577 1 723
2 579 1 723
2 580 1 727
2 581 1 727
2 583 1 730
2 584 1 730
2 585 1 735
2 586 1 735
2 587 1 738
2 588 1 738
2 589 1 741
2 590 1 741
2 591 1 744
2 592 1 744
2 593 1 747
2 595 1 747
2 596 1 750
2 597 1 750
2 598 1 753
2 599 1 753
2 600 1 756
2 601 1 756
2 602 1 759
2 603 1 759
2 604 1 762
2 605 1 762
2 614 1 765
2 615 1 765
2 616 1 768
2 617 1 768
2 618 1 771
2 619 1 771
2 620 1 774
2 621 1 774
2 622 1 777
2 623 1 777
2 624 1 780
2 626 1 780
2 627 1 783
2 628 1 783
2 629 1 786
2 630 1 786
2 631 1 800
2 632 1 800
2 633 1 1034
2 634 1 1034
2 635 1 1037
2 636 1 1037
2 638 1 1037
2 639 1 1037
2 640 1 1042
2 641 1 1042
2 642 1 1042
2 644 1 1042
2 645 1 1042
2 646 1 1042
2 647 1 1042
2 648 1 1042
2 649 1 1042
2 652 1 1042
2 653 1 1053
2 654 1 1053
2 656 1 1053
2 657 1 1053
2 658 1 1053
2 660 1 1053
2 661 1 1053
2 662 1 1053
2 664 1 1053
2 665 1 1053
2 666 1 1070
2 668 1 1070
2 669 1 1070
2 670 1 1070
2 672 1 1075
2 673 1 1075
2 674 1 1075
2 676 1 1075
2 677 1 1075
2 678 1 1075
2 680 1 1075
2 681 1 1075
2 682 1 1075
2 684 1 1075
2 685 1 1086
2 686 1 1086
2 688 1 1086
2 689 1 1086
2 690 1 1086
2 691 1 1086
2 692 1 1086
2 694 1 1086
2 695 1 1086
2 696 1 1086
2 697 1 1102
2 698 1 1102
2 700 1 1102
2 701 1 1102
2 702 1 1102
2 703 1 1102
2 704 1 1102
2 706 1 1102
2 707 1 1102
2 708 1 1102
2 709 1 1113
2 710 1 1113
2 712 1 1113
2 713 1 1113
2 714 1 1113
2 716 1 1113
2 717 1 1113
2 718 1 1113
2 720 1 1113
2 721 1 1113
2 722 1 1129
2 724 1 1129
2 725 1 1129
2 726 1 1133
2 728 1 1133
2 729 1 1133
2 731 1 1137
2 732 1 1137
2 736 1 1146
2 737 1 1146
2 739 1 1146
2 740 1 1146
2 742 1 1146
2 743 1 1146
2 745 1 1146
2 746 1 1146
2 748 1 1146
2 749 1 1146
2 751 1 1157
2 752 1 1157
2 754 1 1157
2 755 1 1157
2 757 1 1157
2 758 1 1157
2 760 1 1157
2 761 1 1157
2 763 1 1157
2 764 1 1157
2 766 1 1173
2 767 1 1173
2 769 1 1173
2 770 1 1173
2 772 1 1178
2 773 1 1178
2 775 1 1178
2 776 1 1178
2 778 1 1178
2 779 1 1190
2 781 1 1190
2 782 1 1190
2 784 1 1190
2 785 1 1195
2 787 1 1195
2 788 1 1195
2 789 1 1195
2 790 1 1200
2 791 1 1200
2 793 1 1200
2 794 1 1200
2 795 1 1205
2 796 1 1205
2 797 1 1205
2 798 1 1205
2 801 1 1216
2 802 1 1216
2 803 1 1219
2 804 1 1219
2 806 1 1222
2 807 1 1222
2 808 1 1225
2 809 1 1225
2 810 1 1228
2 811 1 1228
2 812 1 1231
2 813 1 1231
2 814 1 1234
2 815 1 1234
2 816 1 1237
2 817 1 1237
2 818 1 1240
2 819 1 1240
2 820 1 1243
2 821 1 1243
2 822 1 1246
2 823 1 1246
2 824 1 1251
2 825 1 1251
2 826 1 1254
2 827 1 1254
2 828 1 1257
2 829 1 1257
2 830 1 1260
2 831 1 1260
2 832 1 1263
2 833 1 1263
2 834 1 1266
2 835 1 1266
2 836 1 1496
2 837 1 1496
2 838 1 1499
2 839 1 1499
2 840 1 1502
2 841 1 1502
2 842 1 1502
2 843 1 1506
2 844 1 1506
2 845 1 1506
2 846 1 1510
2 847 1 1510
2 848 1 1513
2 849 1 1513
2 850 1 1516
2 851 1 1516
2 852 1 1553
2 853 1 1553
2 854 1 1553
2 855 1 1557
2 856 1 1557
2 857 1 1557
2 858 1 1561
2 859 1 1561
2 860 1 1578
2 861 1 1578
2 862 1 1582
2 863 1 1582
2 864 1 1585
2 865 1 1585
2 866 1 1588
2 867 1 1588
2 868 1 1591
2 869 1 1591
2 870 1 1591
2 871 1 1591
2 872 1 1596
2 873 1 1596
2 874 1 1596
2 875 1 1600
2 876 1 1600
2 877 1 1600
2 878 1 1600
2 879 1 1600
2 880 1 1606
2 881 1 1606
2 882 1 1606
2 883 1 1606
2 884 1 1606
2 885 1 1612
2 886 1 1612
2 887 1 1615
2 888 1 1615
2 889 1 1615
2 890 1 1619
2 891 1 1619
2 892 1 1619
2 893 1 1619
2 894 1 1624
2 895 1 1624
2 896 1 1624
2 897 1 1628
2 898 1 1628
2 899 1 1631
2 906 1 1631
2 907 1 1634
2 908 1 1634
2 909 1 1637
2 910 1 1637
2 911 1 1637
2 912 1 1637
2 913 1 1642
2 914 1 1642
2 915 1 1642
2 916 1 1642
2 917 1 1647
2 918 1 1647
2 919 1 1647
2 920 1 1651
2 921 1 1651
2 922 1 1651
2 923 1 1651
2 924 1 1656
2 925 1 1656
2 926 1 1656
2 927 1 1676
2 928 1 1676
2 929 1 1676
2 930 1 1676
2 931 1 1681
2 932 1 1681
2 933 1 1681
2 934 1 1681
2 935 1 1686
2 936 1 1686
2 937 1 1686
2 938 1 1690
2 939 1 1690
2 940 1 1708
2 941 1 1708
2 942 1 1770
2 943 1 1770
2 944 1 1773
2 945 1 1773
2 946 1 1778
2 947 1 1778
2 948 1 1781
2 949 1 1781
2 950 1 1795
2 951 1 1795
2 952 1 1798
2 953 1 1798
2 954 1 1801
2 955 1 1801
2 956 1 1804
2 957 1 1804
2 958 1 1824
2 959 1 1824
2 960 1 1827
2 961 1 1827
2 962 1 1833
2 963 1 1833
2 964 1 1836
2 965 1 1836
2 966 1 1836
2 967 1 1836
2 968 1 1841
2 969 1 1841
2 970 1 1841
2 971 1 1841
2 972 1 1841
2 973 1 1841
2 974 1 1848
2 975 1 1848
2 976 1 1848
2 977 1 1852
2 978 1 1852
2 979 1 1852
2 980 1 1856
2 981 1 1856
2 982 1 1856
2 983 1 1856
2 984 1 1856
2 985 1 1856
2 986 1 1863
2 987 1 1863
2 988 1 1863
2 989 1 1863
2 990 1 1863
2 991 1 1863
2 992 1 1870
2 993 1 1870
2 994 1 1870
2 995 1 1870
2 996 1 1875
2 997 1 1875
2 1000 1 1875
2 1001 1 1875
2 1002 1 1880
2 1003 1 1880
2 1004 1 1880
2 1005 1 1880
2 1006 1 1885
2 1007 1 1885
2 1008 1 1888
2 1009 1 1888
2 1010 1 1891
2 1011 1 1891
2 1012 1 1894
2 1013 1 1894
2 1014 1 1897
2 1015 1 1897
2 1016 1 1936
2 1017 1 1936
2 1018 1 1942
2 1019 1 1942
2 1020 1 1945
2 1021 1 1945
2 1022 1 1948
2 1023 1 1948
2 1024 1 1951
2 1025 1 1951
2 1030 1 1954
2 1031 1 1954
2 1035 1 1957
2 1036 1 1957
2 1038 1 1960
2 1039 1 1960
2 1040 1 1963
2 1041 1 1963
2 1043 1 1966
2 1044 1 1966
2 1045 1 2046
2 1046 1 2046
2 1047 1 2049
2 1048 1 2049
2 1049 1 2052
2 1050 1 2052
2 1051 1 2055
2 1052 1 2055
2 1054 1 2058
2 1055 1 2058
2 1056 1 2061
2 1057 1 2061
2 1058 1 2064
2 1059 1 2064
2 1060 1 2067
2 1061 1 2067
2 1062 1 2070
2 1063 1 2070
2 1071 1 2073
2 1072 1 2073
2 1073 1 2076
2 1074 1 2076
2 1076 1 2079
2 1077 1 2079
2 1078 1 2095
2 1079 1 2095
2 1080 1 2098
2 1081 1 2098
2 1082 1 2101
2 1083 1 2101
2 1084 1 2104
2 1085 1 2104
2 1087 1 2107
2 1088 1 2107
2 1089 1 2110
2 1090 1 2110
2 1091 1 2113
2 1092 1 2113
2 1093 1 2113
2 1094 1 2113
2 1095 1 2113
2 1096 1 2120
2 1103 1 2120
2 1104 1 2120
2 1105 1 2120
2 1106 1 2128
2 1107 1 2128
2 1108 1 2128
2 1109 1 2128
2 1110 1 2128
2 1111 1 2128
2 1112 1 2135
2 1114 1 2135
2 1115 1 2135
2 1116 1 2135
2 1117 1 2135
2 1118 1 2141
2 1119 1 2141
2 1120 1 2144
2 1121 1 2144
2 1122 1 2147
2 1123 1 2147
2 1130 1 2150
2 1131 1 2150
2 1132 1 2185
2 1134 1 2185
2 1135 1 2188
2 1136 1 2188
2 1138 1 2191
2 1139 1 2191
2 1147 1 2194
2 1148 1 2194
2 1149 1 2197
2 1150 1 2197
2 1151 1 2201
2 1152 1 2201
2 1153 1 2204
2 1154 1 2204
2 1155 1 2207
2 1156 1 2207
2 1158 1 2210
2 1159 1 2210
2 1160 1 2213
2 1161 1 2213
2 1162 1 2216
2 1163 1 2216
2 1164 1 2219
2 1165 1 2219
2 1166 1 2250
2 1167 1 2250
2 1174 1 2266
2 1175 1 2266
2 1176 1 2269
2 1177 1 2269
2 1179 1 2291
2 1180 1 2291
2 1181 1 2294
2 1182 1 2294
2 1183 1 2359
2 1191 1 2359
2 1192 1 2368
2 1193 1 2368
2 1194 1 2368
2 1196 1 2377
2 1197 1 2377
2 1198 1 2377
2 1199 1 2377
2 1201 1 2382
2 1202 1 2382
2 1203 1 2382
2 1204 1 2391
2 1206 1 2391
2 1207 1 2391
2 1208 1 2395
2 1209 1 2395
2 1217 1 2395
2 1218 1 2395
2 1220 1 2417
2 1221 1 2417
2 1223 1 2417
2 1224 1 2421
2 1226 1 2421
2 1227 1 2421
2 1229 1 2425
2 1230 1 2425
2 1232 1 2434
2 1233 1 2434
2 1235 1 2437
2 1236 1 2437
2 1238 1 2440
2 1239 1 2440
2 1241 1 2443
2 1242 1 2443
2 1244 1 2446
2 1245 1 2446
2 1247 1 2449
2 1248 1 2449
2 1252 1 2454
2 1253 1 2454
2 1255 1 2457
2 1256 1 2457
2 1258 1 2460
2 1259 1 2460
2 1261 1 2463
2 1262 1 2463
2 1264 1 2466
2 1265 1 2466
2 1267 1 2469
2 1268 1 2469
2 1270 1 2472
2 1271 1 2472
2 1272 1 2475
2 1273 1 2475
2 1274 1 2478
2 1278 1 2478
2 1279 1 2481
2 1280 1 2481
2 1281 1 2484
2 1282 1 2484
2 1283 1 2487
2 1284 1 2487
2 1285 1 2490
2 1286 1 2490
2 1287 1 2493
2 1288 1 2493
2 1289 1 2521
2 1290 1 2521
2 1291 1 2531
2 1292 1 2531
2 1293 1 2534
2 1294 1 2534
2 1295 1 2537
2 1296 1 2537
2 1297 1 2540
2 1298 1 2540
2 1299 1 2603
2 1300 1 2603
2 1301 1 2603
2 1303 1 2613
2 1304 1 2613
2 1305 1 2613
2 1306 1 2621
2 1307 1 2621
2 1308 1 2624
2 1309 1 2624
2 1310 1 2624
2 1311 1 2638
2 1312 1 2638
2 1313 1 2638
2 1314 1 2638
2 1315 1 2646
2 1316 1 2646
2 1317 1 2646
2 1318 1 2646
2 1319 1 2659
2 1320 1 2659
2 1321 1 2659
2 1322 1 2681
2 1323 1 2681
2 1324 1 2684
2 1325 1 2684
2 1326 1 2687
2 1327 1 2687
2 1328 1 2690
2 1329 1 2690
2 1330 1 2703
2 1331 1 2703
2 1332 1 2729
2 1333 1 2729
2 1334 1 2729
2 1335 1 2729
2 1336 1 2738
2 1337 1 2738
2 1338 1 2738
2 1339 1 2738
2 1340 1 2761
2 1341 1 2761
2 1342 1 2761
2 1343 1 2761
2 1344 1 2766
2 1345 1 2766
2 1346 1 2766
2 1347 1 2766
2 1348 1 2793
2 1349 1 2793
2 1350 1 2796
2 1356 1 2796
2 1357 1 2796
2 1358 1 2800
2 1359 1 2800
2 1360 1 2803
2 1361 1 2803
2 1362 1 2806
2 1363 1 2806
2 1364 1 2817
2 1365 1 2817
2 1366 1 2820
2 1367 1 2820
2 1368 1 2820
2 1369 1 2820
2 1370 1 2820
2 1371 1 2826
2 1372 1 2826
2 1373 1 2831
2 1374 1 2831
2 1375 1 2831
2 1376 1 2831
2 1377 1 2831
2 1378 1 2841
2 1379 1 2841
2 1380 1 2844
2 1381 1 2844
2 1382 1 2844
2 1383 1 2844
2 1384 1 2844
2 1385 1 2854
2 1386 1 2854
2 1387 1 2854
2 1388 1 2854
2 1389 1 2859
2 1390 1 2859
2 1391 1 2859
2 1392 1 2859
2 1393 1 2859
2 1394 1 2869
2 1400 1 2869
2 1401 1 2869
2 1402 1 2869
2 1403 1 2874
2 1404 1 2874
2 1405 1 2877
2 1406 1 2877
2 1407 1 2882
2 1408 1 2882
2 1409 1 2885
2 1410 1 2885
2 1411 1 2888
2 1412 1 2888
2 1413 1 2931
2 1414 1 2931
2 1415 1 2972
2 1416 1 2972
2 1417 1 2975
2 1418 1 2975
2 1419 1 2978
2 1420 1 2978
2 1421 1 2981
2 1428 1 2981
2 1429 1 2986
2 1430 1 2986
2 1431 1 2989
2 1432 1 2989
2 1433 1 2992
2 1434 1 2992
2 1435 1 2995
2 1436 1 2995
2 1437 1 2998
2 1438 1 2998
2 1439 1 3001
2 1442 1 3001
2 1443 1 3004
2 1444 1 3004
2 1445 1 3010
2 1446 1 3010
2 1447 1 3013
2 1497 1 3013
2 1498 1 3016
2 1500 1 3016
2 1501 1 3019
2 1503 1 3019
2 1504 1 3022
2 1505 1 3022
2 1507 1 3025
2 1508 1 3025
2 1509 1 3030
2 1511 1 3030
2 1512 1 3030
2 1514 1 3030
2 1515 1 3039
2 1517 1 3039
2 1518 1 3039
2 1554 1 3039
2 1555 1 3050
2 1556 1 3050
2 1558 1 3061
2 1559 1 3061
2 1560 1 3076
2 1562 1 3076
2 1563 1 3088
2 1579 1 3088
2 1580 1 3091
2 1583 1 3091
2 1584 1 3110
2 1586 1 3110
2 1587 1 3113
2 1589 1 3113
2 1590 1 3137
2 1592 1 3137
2 1593 1 3140
2 1594 1 3140
2 1595 1 3143
2 1597 1 3143
2 1598 1 3146
2 1599 1 3146
2 1601 1 3149
2 1602 1 3149
2 1603 1 3152
2 1604 1 3152
2 1605 1 3157
2 1607 1 3157
2 1608 1 3160
2 1609 1 3160
2 1610 1 3163
2 1611 1 3163
2 1613 1 3166
2 1614 1 3166
2 1616 1 3169
2 1617 1 3169
2 1618 1 3172
2 1620 1 3172
2 1621 1 3180
2 1622 1 3180
2 1623 1 3238
2 1625 1 3238
2 1626 1 3241
2 1627 1 3241
2 1629 1 3244
2 1630 1 3244
2 1632 1 3247
2 1633 1 3247
2 1635 1 3250
2 1636 1 3250
2 1638 1 3253
2 1639 1 3253
2 1640 1 3256
2 1641 1 3256
2 1643 1 3259
2 1644 1 3259
2 1645 1 3262
2 1646 1 3262
2 1648 1 3265
2 1649 1 3265
2 1650 1 3268
2 1652 1 3268
2 1653 1 3271
2 1654 1 3271
2 1655 1 3274
2 1657 1 3274
2 1658 1 3277
2 1659 1 3277
2 1660 1 3315
2 1661 1 3315
2 1662 1 3318
2 1663 1 3318
2 1664 1 3321
2 1665 1 3321
2 1666 1 3324
2 1667 1 3324
2 1668 1 3327
2 1669 1 3327
2 1670 1 3330
2 1671 1 3330
2 1672 1 3340
2 1673 1 3340
2 1674 1 3344
2 1675 1 3344
2 1677 1 3348
2 1678 1 3348
2 1679 1 3352
2 1680 1 3352
2 1682 1 3356
2 1683 1 3356
2 1684 1 3360
2 1685 1 3360
2 1687 1 3364
2 1688 1 3364
2 1689 1 3367
2 1691 1 3367
2 1692 1 3370
2 1693 1 3370
2 1694 1 3374
2 1695 1 3374
2 1696 1 3378
2 1697 1 3378
2 1698 1 3382
2 1699 1 3382
2 1700 1 3386
2 1701 1 3386
2 1702 1 3390
2 1703 1 3390
2 1704 1 3394
2 1705 1 3394
2 1706 1 3397
2 1707 1 3397
2 1709 1 3450
2 1710 1 3450
2 1711 1 3453
2 1712 1 3453
2 1713 1 3456
2 1714 1 3456
2 1715 1 3459
2 1716 1 3459
2 1717 1 3522
2 1718 1 3522
2 1719 1 3525
2 1720 1 3525
2 1721 1 3528
2 1722 1 3528
2 1723 1 3531
2 1724 1 3531
2 1725 1 3534
2 1727 1 3534
2 1728 1 3537
2 1729 1 3537
2 1730 1 3540
2 1731 1 3540
2 1732 1 3543
2 1733 1 3543
2 1734 1 3576
2 1735 1 3576
2 1736 1 3579
2 1737 1 3579
2 1738 1 3585
2 1739 1 3585
2 1740 1 3588
2 1741 1 3588
2 1742 1 3600
2 1743 1 3600
2 1744 1 3603
2 1745 1 3603
2 1746 1 3603
2 1747 1 3603
2 1748 1 3608
2 1749 1 3608
2 1750 1 3608
2 1751 1 3612
2 1752 1 3612
2 1753 1 3616
2 1754 1 3616
2 1755 1 3616
2 1756 1 3616
2 1757 1 3616
2 1758 1 3622
2 1759 1 3622
2 1760 1 3622
2 1761 1 3622
2 1762 1 3635
2 1763 1 3635
2 1764 1 3635
2 1765 1 3635
2 1766 1 3640
2 1767 1 3640
2 1768 1 3640
2 1769 1 3644
2 1771 1 3644
2 1772 1 3648
2 1774 1 3648
2 1775 1 3648
2 1779 1 3648
2 1780 1 3648
2 1782 1 3654
2 1783 1 3654
2 1786 1 3654
2 1787 1 3654
2 1788 1 3723
2 1789 1 3723
2 1790 1 3737
2 1791 1 3737
2 1792 1 3754
2 1793 1 3754
2 1794 1 3754
2 1796 1 3758
2 1797 1 3758
2 1799 1 3762
2 1800 1 3762
2 1802 1 3767
2 1803 1 3767
2 1805 1 3767
2 1806 1 3771
2 1812 1 3771
2 1825 1 3775
2 1826 1 3775
2 1828 1 3780
2 1829 1 3780
2 1834 1 3790
2 1835 1 3790
2 1837 1 3823
2 1838 1 3823
2 1839 1 3827
2 1840 1 3827
2 1842 1 3840
2 1843 1 3840
2 1844 1 3843
2 1845 1 3843
2 1846 1 3843
2 1847 1 3852
2 1849 1 3852
2 1850 1 3859
2 1851 1 3859
2 1853 1 3864
2 1854 1 3864
2 1855 1 3870
2 1857 1 3870
2 1858 1 3877
2 1859 1 3877
