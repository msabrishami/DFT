1 0 0 5 0
1 1 0 2 0
1 2 0 3 0
1 3 0 5 0
1 4 0 1 0
1 5 0 3 0
1 6 0 4 0
1 7 0 4 0
1 8 0 2 0
1 9 0 3 0
1 10 0 4 0
1 11 0 1 0
1 12 0 1 0
1 13 0 1 0
1 14 0 1 0
1 15 0 2 0
1 16 0 2 0
1 17 0 1 0
1 18 0 1 0
1 19 0 1 0
1 20 0 1 0
1 21 0 1 0
1 22 0 1 0
1 23 0 3 0
1 24 0 3 0
1 25 0 1 0
1 26 0 2 0
1 27 0 2 0
1 28 0 4 0
1 29 0 4 0
1 30 0 3 0
1 31 0 5 0
1 32 0 3 0
1 33 0 2 0
1 34 0 2 0
1 35 0 2 0
1 36 0 2 0
1 37 0 1 0
1 38 0 2 0
1 39 0 1 0
1 40 0 3 0
1 41 0 4 0
1 42 0 5 0
1 43 0 4 0
1 44 0 4 0
1 45 0 4 0
1 46 0 5 0
1 47 0 5 0
1 48 0 3 0
1 49 0 4 0
1 50 0 8 0
1 51 0 3 0
1 52 0 8 0
1 53 0 6 0
1 54 0 3 0
1 55 0 1 0
1 56 0 1 0
1 57 0 3 0
1 58 0 1 0
1 59 0 2 0
0 60 7 1 2 13 12
0 61 5 4 1 25
0 62 3 2 2 19 20
3 63 7 0 2 18 17
0 64 5 1 1 4
2 65 1 0 
2 66 1 0 
2 67 1 0 
2 68 1 0 
2 69 1 0 
2 70 1 1 
2 71 1 1 
2 72 1 2 
2 73 1 2 
2 74 1 2 
2 75 1 3 
2 76 1 3 
2 77 1 3 
2 78 1 3 
2 79 1 3 
2 80 1 5 
2 81 1 5 
2 82 1 5 
2 83 1 6 
2 84 1 6 
2 85 1 6 
2 86 1 6 
2 87 1 7 
2 88 1 7 
2 89 1 7 
2 90 1 7 
2 91 1 8 
2 92 1 8 
2 93 1 9 
2 94 1 9 
2 95 1 9 
2 96 1 10 
2 97 1 10 
2 98 1 10 
2 99 1 10 
2 100 1 15 
2 101 1 15 
2 102 1 16 
2 103 1 16 
2 104 1 23 
2 105 1 23 
2 106 1 23 
2 107 1 24 
2 108 1 24 
2 109 1 24 
2 110 1 26 
2 111 1 26 
2 112 1 27 
2 113 1 27 
2 114 1 28 
2 115 1 28 
2 116 1 28 
2 117 1 28 
2 118 1 29 
2 119 1 29 
2 120 1 29 
2 121 1 29 
2 122 1 30 
2 123 1 30 
2 124 1 30 
2 125 1 31 
2 126 1 31 
2 127 1 31 
2 128 1 31 
2 129 1 31 
2 130 1 32 
2 131 1 32 
2 132 1 32 
2 133 1 33 
2 134 1 33 
2 135 1 34 
2 136 1 34 
2 137 1 35 
2 138 1 35 
2 139 1 36 
2 140 1 36 
2 141 1 38 
2 142 1 38 
2 143 1 40 
2 144 1 40 
2 145 1 40 
2 146 1 41 
2 147 1 41 
2 148 1 41 
2 149 1 41 
2 150 1 42 
2 151 1 42 
2 152 1 42 
2 153 1 42 
2 154 1 42 
2 155 1 43 
2 156 1 43 
2 157 1 43 
2 158 1 43 
2 159 1 44 
2 160 1 44 
2 161 1 44 
2 162 1 44 
2 163 1 45 
2 164 1 45 
2 165 1 45 
2 166 1 45 
2 167 1 46 
2 168 1 46 
2 169 1 46 
2 170 1 46 
2 171 1 46 
2 172 1 47 
2 173 1 47 
2 174 1 47 
2 175 1 47 
2 176 1 47 
2 177 1 48 
2 178 1 48 
2 179 1 48 
2 180 1 49 
2 181 1 49 
2 182 1 49 
2 183 1 49 
2 184 1 50 
2 185 1 50 
2 186 1 50 
2 187 1 50 
2 188 1 50 
2 189 1 50 
2 190 1 50 
2 191 1 50 
2 192 1 51 
2 193 1 51 
2 194 1 51 
2 195 1 52 
2 196 1 52 
2 197 1 52 
2 198 1 52 
2 199 1 52 
2 200 1 52 
2 201 1 52 
2 202 1 52 
2 203 1 53 
2 204 1 53 
2 205 1 53 
2 206 1 53 
2 207 1 53 
2 208 1 53 
2 209 1 54 
2 210 1 54 
2 211 1 54 
2 212 1 57 
2 213 1 57 
2 214 1 57 
2 215 1 59 
2 216 1 59 
0 217 7 1 2 180 215
0 218 5 1 1 139
0 219 5 1 1 137
0 220 5 1 1 135
0 221 5 3 1 133
0 222 5 1 1 141
0 223 7 1 2 37 134
0 224 6 1 2 114 181
0 225 6 1 2 56 209
0 226 6 1 2 55 210
0 227 5 2 1 189
0 228 5 5 1 182
0 229 5 1 1 213
0 230 6 1 2 87 96
0 231 5 3 1 208
0 232 6 1 2 118 183
0 233 6 1 2 58 211
0 234 5 6 1 194
0 235 7 3 2 39 97
0 236 5 2 1 91
0 237 5 3 1 77
0 238 5 3 1 144
0 239 5 2 1 149
0 240 5 3 1 153
0 241 5 4 1 158
0 242 5 4 1 161
0 243 5 4 1 166
0 244 5 3 1 171
0 245 5 3 1 175
0 246 5 2 1 179
0 247 5 3 1 121
0 248 5 3 1 110
0 249 5 3 1 113
0 250 5 3 1 116
0 251 5 2 1 129
0 252 5 4 1 105
0 253 5 4 1 109
0 254 5 3 1 123
0 255 5 2 1 132
0 256 6 1 2 67 95
0 257 5 3 1 70
0 258 7 1 2 11 72
0 259 5 4 1 98
0 260 5 2 1 102
0 261 5 2 1 100
0 262 7 1 2 73 78
0 263 6 1 2 71 74
0 264 6 1 2 68 79
0 265 5 3 1 80
0 266 6 1 2 81 103
0 267 5 1 1 86
0 268 6 1 2 82 101
0 269 5 4 1 90
0 270 5 1 1 69
2 271 1 61 
2 272 1 61 
2 273 1 61 
2 274 1 61 
2 275 1 62 
2 276 1 62 
0 277 6 1 2 225 224
0 278 6 1 2 233 232
3 279 7 0 2 21 275
3 280 7 0 2 22 276
3 281 4 0 2 264 263
3 282 4 0 2 267 266
0 283 4 2 2 270 64
2 284 1 221 
2 285 1 221 
2 286 1 221 
2 287 1 227 
2 288 1 227 
2 289 1 228 
2 290 1 228 
2 291 1 228 
2 292 1 228 
2 293 1 228 
2 294 1 231 
2 295 1 231 
2 296 1 231 
2 297 1 234 
2 298 1 234 
2 299 1 234 
2 300 1 234 
2 301 1 234 
2 302 1 234 
2 303 1 235 
2 304 1 235 
2 305 1 235 
2 306 1 236 
2 307 1 236 
2 308 1 237 
2 309 1 237 
2 310 1 237 
2 311 1 238 
2 312 1 238 
2 313 1 238 
2 314 1 239 
2 315 1 239 
2 316 1 240 
2 317 1 240 
2 318 1 240 
2 319 1 241 
2 320 1 241 
2 321 1 241 
2 322 1 241 
2 323 1 242 
2 324 1 242 
2 325 1 242 
2 326 1 242 
2 327 1 243 
2 328 1 243 
2 329 1 243 
2 330 1 243 
2 331 1 244 
2 332 1 244 
2 333 1 244 
2 334 1 245 
2 335 1 245 
2 336 1 245 
2 337 1 246 
2 338 1 246 
2 339 1 247 
2 340 1 247 
2 341 1 247 
2 342 1 248 
2 343 1 248 
2 344 1 248 
2 345 1 249 
2 346 1 249 
2 347 1 249 
2 348 1 250 
2 349 1 250 
2 350 1 250 
2 351 1 251 
2 352 1 251 
2 353 1 252 
2 354 1 252 
2 355 1 252 
2 356 1 252 
2 357 1 253 
2 358 1 253 
2 359 1 253 
2 360 1 253 
2 361 1 254 
2 362 1 254 
2 363 1 254 
2 364 1 255 
2 365 1 255 
2 366 1 257 
2 367 1 257 
2 368 1 257 
2 369 1 259 
2 370 1 259 
2 371 1 259 
2 372 1 259 
2 373 1 260 
2 374 1 260 
2 375 1 261 
2 376 1 261 
2 377 1 265 
2 378 1 265 
2 379 1 265 
2 380 1 269 
2 381 1 269 
2 382 1 269 
2 383 1 269 
0 384 4 1 2 289 357
0 385 4 1 2 290 353
0 386 4 1 2 284 308
0 387 4 1 2 285 306
0 388 4 1 2 286 366
0 389 4 1 2 291 272
0 390 4 1 2 292 345
0 391 4 1 2 293 343
0 392 4 1 2 88 309
0 393 4 1 2 76 380
0 394 4 1 2 369 375
0 395 4 1 2 310 367
0 396 4 1 2 216 377
0 397 6 1 2 177 335
0 398 6 1 2 174 337
0 399 6 1 2 148 313
0 400 6 1 2 145 315
0 401 6 1 2 164 325
0 402 6 1 2 160 329
0 403 4 1 2 156 317
0 404 4 1 2 152 321
0 405 6 1 2 157 318
0 406 6 1 2 154 322
0 407 4 1 2 165 326
0 408 4 1 2 162 330
0 409 4 1 2 178 336
0 410 4 1 2 176 338
0 411 6 1 2 130 362
0 412 6 1 2 122 364
0 413 6 1 2 112 344
0 414 6 1 2 111 347
0 415 6 1 2 107 355
0 416 6 1 2 104 359
0 417 4 1 2 127 349
0 418 4 1 2 115 351
0 419 6 1 2 128 350
0 420 6 1 2 117 352
0 421 4 1 2 108 356
0 422 4 1 2 106 360
0 423 4 1 2 131 363
0 424 4 1 2 124 365
0 425 4 1 2 256 368
0 426 4 1 2 371 381
0 427 4 1 2 372 373
0 428 4 2 2 374 376
0 429 4 1 2 379 382
3 430 4 0 2 268 383
2 431 1 283 
2 432 1 283 
0 433 4 1 2 393 392
0 434 6 1 2 394 89
0 435 6 1 2 398 397
0 436 6 2 2 400 399
0 437 6 1 2 402 401
0 438 4 1 2 404 403
0 439 6 1 2 406 405
0 440 4 1 2 408 407
0 441 4 1 2 410 409
0 442 6 1 2 412 411
0 443 6 2 2 414 413
0 444 6 1 2 416 415
0 445 4 1 2 418 417
0 446 6 1 2 420 419
0 447 4 1 2 422 421
0 448 4 1 2 424 423
0 449 6 3 2 258 425
3 450 6 0 2 426 83
3 451 6 0 2 427 84
0 452 7 2 2 262 431
0 453 6 2 2 429 85
0 454 6 4 2 92 432
2 455 1 428 
2 456 1 428 
0 457 6 1 2 434 66
0 458 6 2 2 396 455
0 459 6 1 2 438 437
0 460 6 1 2 440 439
0 461 6 2 2 445 444
0 462 6 2 2 447 446
3 463 6 0 2 99 456
2 464 1 436 
2 465 1 436 
2 466 1 443 
2 467 1 443 
2 468 1 449 
2 469 1 449 
2 470 1 449 
2 471 1 452 
2 472 1 452 
2 473 1 453 
2 474 1 453 
2 475 1 454 
2 476 1 454 
2 477 1 454 
2 478 1 454 
0 479 4 1 2 303 475
0 480 4 1 2 230 468
0 481 4 1 2 433 476
0 482 4 1 2 457 307
0 483 6 2 2 460 459
0 484 4 2 2 273 466
0 485 7 2 2 274 467
0 486 4 1 2 469 370
3 487 4 0 2 470 378
3 488 6 0 2 472 473
3 489 5 0 1 474
3 490 5 0 1 478
2 491 1 458 
2 492 1 458 
2 493 1 461 
2 494 1 461 
2 495 1 462 
2 496 1 462 
0 497 6 4 2 479 93
0 498 6 4 2 60 480
0 499 6 2 2 490 75
0 500 6 1 2 481 305
0 501 6 1 2 395 482
0 502 4 1 2 492 477
0 503 6 1 2 493 495
0 504 7 1 2 494 496
3 505 7 0 2 486 14
3 506 6 0 2 489 471
2 507 1 483 
2 508 1 483 
2 509 1 484 
2 510 1 484 
2 511 1 485 
2 512 1 485 
0 513 7 8 2 501 500
0 514 7 4 2 502 94
0 515 6 1 2 125 507
0 516 3 1 2 126 508
0 517 4 1 2 509 511
0 518 3 1 2 510 512
2 519 1 497 
2 520 1 497 
2 521 1 497 
2 522 1 497 
2 523 1 498 
2 524 1 498 
2 525 1 498 
2 526 1 498 
2 527 1 499 
2 528 1 499 
0 529 4 1 2 523 316
0 530 4 1 2 218 519
0 531 4 1 2 219 520
0 532 4 1 2 220 521
0 533 4 1 2 222 522
0 534 4 4 2 527 491
0 535 4 1 2 525 331
0 536 5 5 1 526
0 537 3 1 2 528 304
0 538 7 2 2 516 515
0 539 6 1 2 517 503
0 540 6 1 2 504 518
2 541 1 513 
2 542 1 513 
2 543 1 513 
2 544 1 513 
2 545 1 513 
2 546 1 513 
2 547 1 513 
2 548 1 513 
2 549 1 514 
2 550 1 514 
2 551 1 514 
2 552 1 514 
0 553 4 1 2 541 271
0 554 4 1 2 542 358
0 555 4 1 2 543 354
0 556 4 1 2 544 342
0 557 4 1 2 545 339
0 558 4 1 2 546 348
0 559 4 1 2 547 346
0 560 6 4 2 537 65
0 561 4 1 2 548 361
0 562 6 3 2 540 539
2 563 1 534 
2 564 1 534 
2 565 1 534 
2 566 1 534 
2 567 1 536 
2 568 1 536 
2 569 1 536 
2 570 1 536 
2 571 1 536 
2 572 1 538 
2 573 1 538 
0 574 6 1 2 143 567
0 575 4 1 2 530 563
0 576 4 1 2 553 386
0 577 4 1 2 531 564
0 578 4 1 2 554 387
0 579 4 1 2 532 565
0 580 4 1 2 555 388
0 581 4 1 2 533 566
0 582 4 1 2 556 223
0 583 6 1 2 155 568
0 584 4 1 2 557 549
0 585 4 1 2 558 550
0 586 4 1 2 559 551
0 587 6 1 2 159 570
0 588 6 1 2 172 571
0 589 4 1 2 561 552
0 590 6 1 2 464 572
0 591 3 1 2 465 573
2 592 1 560 
2 593 1 560 
2 594 1 560 
2 595 1 560 
2 596 1 562 
2 597 1 562 
2 598 1 562 
0 599 6 3 2 576 575
0 600 6 3 2 578 577
0 601 6 2 2 580 579
0 602 6 2 2 582 581
0 603 6 1 2 140 592
0 604 6 1 2 138 593
0 605 6 1 2 136 594
0 606 6 1 2 142 595
0 607 6 3 2 591 590
0 608 6 1 2 119 596
0 609 4 1 2 120 597
0 610 5 2 1 598
0 611 6 3 2 584 603
0 612 6 3 2 585 604
0 613 6 2 2 586 605
0 614 6 2 2 589 606
2 615 1 599 
2 616 1 599 
2 617 1 599 
2 618 1 600 
2 619 1 600 
2 620 1 600 
2 621 1 601 
2 622 1 601 
2 623 1 602 
2 624 1 602 
2 625 1 607 
2 626 1 607 
2 627 1 607 
2 628 1 610 
2 629 1 610 
0 630 6 1 2 203 615
0 631 6 1 2 196 618
0 632 6 1 2 204 621
0 633 5 2 1 619
0 634 6 3 2 150 616
0 635 4 4 2 151 617
0 636 6 2 2 147 620
0 637 5 2 1 622
0 638 5 2 1 623
0 639 6 1 2 205 624
0 640 6 1 2 625 332
0 641 5 2 1 626
0 642 4 1 2 627 333
0 643 6 1 2 340 628
0 644 4 1 2 341 629
2 645 1 611 
2 646 1 611 
2 647 1 611 
2 648 1 612 
2 649 1 612 
2 650 1 612 
2 651 1 613 
2 652 1 613 
2 653 1 614 
2 654 1 614 
0 655 6 1 2 631 524
0 656 6 1 2 574 632
0 657 6 1 2 583 639
0 658 6 1 2 206 645
0 659 7 1 2 200 648
0 660 5 2 1 649
0 661 4 3 2 167 646
0 662 6 3 2 168 647
0 663 6 2 2 163 650
0 664 5 2 1 651
0 665 6 1 2 207 652
0 666 4 3 2 173 653
0 667 5 2 1 654
0 668 6 1 2 643 608
0 669 4 1 2 644 609
2 670 1 633 
2 671 1 633 
2 672 1 634 
2 673 1 634 
2 674 1 634 
2 675 1 635 
2 676 1 635 
2 677 1 635 
2 678 1 635 
2 679 1 636 
2 680 1 636 
2 681 1 637 
2 682 1 637 
2 683 1 638 
2 684 1 638 
2 685 1 641 
2 686 1 641 
0 687 4 1 2 676 297
0 688 5 3 1 673
0 689 6 1 2 655 146
0 690 4 1 2 670 294
0 691 4 1 2 217 656
0 692 6 2 2 671 314
0 693 6 2 2 681 311
0 694 4 2 2 682 312
0 695 6 3 2 683 319
0 696 4 2 2 684 320
0 697 4 1 2 389 657
0 698 4 1 2 659 569
0 699 6 1 2 587 665
0 700 6 1 2 169 685
0 701 4 1 2 170 686
0 702 6 1 2 442 668
0 703 6 1 2 448 669
2 704 1 660 
2 705 1 660 
2 706 1 661 
2 707 1 661 
2 708 1 661 
2 709 1 662 
2 710 1 662 
2 711 1 662 
2 712 1 663 
2 713 1 663 
2 714 1 664 
2 715 1 664 
2 716 1 666 
2 717 1 666 
2 718 1 666 
2 719 1 667 
2 720 1 667 
0 721 6 1 2 687 672
0 722 4 1 2 690 385
0 723 5 2 1 710
0 724 4 1 2 704 295
0 725 4 1 2 698 327
0 726 6 2 2 705 328
0 727 6 2 2 714 323
0 728 4 2 2 715 324
0 729 4 1 2 391 699
0 730 5 2 1 716
0 731 4 1 2 296 719
0 732 4 1 2 302 718
0 733 4 3 2 720 334
0 734 6 1 2 640 700
0 735 4 1 2 642 701
3 736 6 0 2 703 702
2 737 1 688 
2 738 1 688 
2 739 1 688 
2 740 1 692 
2 741 1 692 
2 742 1 693 
2 743 1 693 
2 744 1 694 
2 745 1 694 
2 746 1 695 
2 747 1 695 
2 748 1 695 
2 749 1 696 
2 750 1 696 
0 751 4 1 2 737 675
0 752 6 1 2 195 739
0 753 6 2 2 740 679
0 754 6 1 2 197 744
0 755 5 2 1 745
0 756 6 1 2 198 749
0 757 5 3 1 750
0 758 4 1 2 724 390
0 759 6 1 2 435 734
0 760 6 1 2 441 735
2 761 1 723 
2 762 1 723 
2 763 1 726 
2 764 1 726 
2 765 1 727 
2 766 1 727 
2 767 1 728 
2 768 1 728 
2 769 1 730 
2 770 1 730 
2 771 1 733 
2 772 1 733 
2 773 1 733 
0 774 6 1 2 752 721
0 775 4 1 2 761 707
0 776 6 1 2 199 762
0 777 6 1 2 758 226
0 778 7 3 2 763 712
0 779 6 1 2 212 769
0 780 6 1 2 201 767
0 781 5 2 1 768
0 782 4 1 2 717 771
0 783 5 3 1 772
0 784 6 1 2 202 773
3 785 6 0 2 760 759
2 786 1 753 
2 787 1 753 
2 788 1 755 
2 789 1 755 
2 790 1 757 
2 791 1 757 
2 792 1 757 
0 793 4 1 2 384 774
0 794 5 2 1 786
0 795 4 1 2 787 298
0 796 6 2 2 742 788
0 797 3 1 2 677 791
0 798 6 3 2 748 792
0 799 4 1 2 782 214
2 800 1 778 
2 801 1 778 
2 802 1 778 
2 803 1 781 
2 804 1 781 
2 805 1 783 
2 806 1 783 
2 807 1 783 
0 808 6 1 2 193 800
0 809 6 2 2 779 805
0 810 6 3 2 766 804
0 811 6 1 2 770 806
0 812 6 1 2 732 807
2 813 1 794 
2 814 1 794 
2 815 1 796 
2 816 1 796 
2 817 1 798 
2 818 1 798 
2 819 1 798 
0 820 5 2 1 815
0 821 4 1 2 816 299
0 822 4 1 2 819 300
0 823 4 1 2 229 811
0 824 6 1 2 784 812
2 825 1 809 
2 826 1 809 
2 827 1 810 
2 828 1 810 
2 829 1 810 
0 830 7 2 2 775 825
0 831 5 2 1 826
0 832 4 1 2 829 301
0 833 4 1 2 799 823
0 834 4 1 2 824 278
2 835 1 820 
2 836 1 820 
0 837 6 1 2 833 191
2 838 1 830 
2 839 1 830 
2 840 1 831 
2 841 1 831 
0 842 4 1 2 838 840
0 843 4 1 2 839 287
0 844 3 1 2 708 841
0 845 6 1 2 588 837
0 846 6 1 2 842 188
0 847 4 1 2 843 192
0 848 6 3 2 844 711
0 849 4 1 2 731 845
0 850 6 1 2 658 846
0 851 4 1 2 847 706
3 852 6 0 2 834 849
2 853 1 848 
2 854 1 848 
2 855 1 848 
0 856 4 1 2 535 850
0 857 6 1 2 851 709
0 858 6 1 2 801 853
0 859 3 1 2 802 854
0 860 6 1 2 764 855
0 861 6 1 2 776 857
0 862 6 1 2 859 858
0 863 6 2 2 860 713
0 864 4 1 2 861 277
0 865 4 1 2 862 288
2 866 1 863 
2 867 1 863 
0 868 6 1 2 866 765
3 869 6 0 2 864 856
0 870 4 1 2 725 865
0 871 5 2 1 867
0 872 6 2 2 868 803
0 873 6 1 2 870 808
2 874 1 871 
2 875 1 871 
3 876 3 0 2 873 777
0 877 4 1 2 874 827
0 878 7 1 2 875 828
2 879 1 872 
2 880 1 872 
0 881 6 1 2 879 746
0 882 5 3 1 880
0 883 4 1 2 878 877
0 884 6 1 2 881 790
0 885 6 1 2 883 190
2 886 1 882 
2 887 1 882 
2 888 1 882 
0 889 4 1 2 751 884
0 890 4 1 2 678 886
0 891 4 1 2 887 817
0 892 7 1 2 888 818
0 893 6 1 2 780 885
0 894 6 1 2 890 747
0 895 4 1 2 892 891
0 896 4 1 2 832 893
0 897 7 2 2 894 797
0 898 6 1 2 895 187
3 899 6 0 2 729 896
0 900 6 1 2 756 898
2 901 1 897 
2 902 1 897 
0 903 4 1 2 738 901
0 904 6 3 2 674 902
0 905 4 1 2 822 900
0 906 4 1 2 903 889
3 907 6 0 2 697 905
2 908 1 904 
2 909 1 904 
2 910 1 904 
0 911 6 1 2 906 184
0 912 4 1 2 813 908
0 913 7 1 2 814 909
0 914 6 1 2 741 910
0 915 6 1 2 630 911
0 916 4 1 2 913 912
0 917 6 3 2 914 680
0 918 4 1 2 529 915
0 919 6 1 2 916 185
2 920 1 917 
2 921 1 917 
2 922 1 917 
3 923 6 0 2 793 918
0 924 6 1 2 689 919
0 925 4 1 2 835 920
0 926 7 1 2 836 921
0 927 6 1 2 922 743
0 928 4 1 2 795 924
0 929 4 1 2 926 925
3 930 6 0 2 927 789
3 931 6 0 2 722 928
0 932 6 1 2 929 186
0 933 6 1 2 754 932
0 934 4 1 2 821 933
3 935 6 0 2 691 934
