1 1 0 1 0 
1 2 0 1 0 
1 3 0 1 0 
0 4 7 4 1 1 
2 5 1 4 
2 6 1 4 
2 7 1 4 
2 8 1 4 
0 9 7 2 1 2 
2 10 1 9 
2 11 1 9 
0 12 7 2 1 3 
2 13 1 12 
2 14 1 12 
0 15 5 2 1 8 
2 16 1 15 
2 17 1 15 
0 18 5 1 1 10 
0 19 5 1 1 14 
0 20 7 2 2 18 13 
2 21 1 20 
2 22 1 20 
0 23 7 3 2 11 19 
2 24 1 23 
2 25 1 23 
2 26 1 23 
0 27 7 1 2 16 21 
0 28 3 2 2 22 24 
2 29 1 28 
2 30 1 28 
0 31 7 1 2 26 17 
0 32 5 2 1 30 
2 33 1 32 
2 34 1 32 
0 35 7 1 2 7 33 
0 36 3 1 2 34 25 
0 37 7 1 2 6 36 
3 38 3 0 2 37 27 
3 39 7 0 2 5 29 
3 40 3 0 2 35 31 
