1 1	0 1	0	
1 2	0 1	0	
1 3	0 2	0	
2 8	1 3	
2 9	1 3	
1 4	0 2	0	
2 10 1 4		
2 11 1 4		
1 5	0 2	0	
2 12 1 5		
2 13 1 5		
1 6	0 1	0	
1 7	0 1	0	
0 14 7 1 2 1 2
0 15 7 1 2 8 10
0 16 5 1 1 9
0 17 5 1 1 11
0 18 5 1 1 13
0 19 7 1 3 12 6 7
0 20 3 1 2 14 15
0 21 3 1 3 16 17 18
3 22 7 0 3 20 21 19