2	8192	1	103			
3	1	0	0	0	
2	8194	1	106			
2	8195	1	106			
1	4	0	7	0	
2	8193	1	103			
2	8198	1	123			
2	8196	1	109			
2	8197	1	109			
2	8199	1	123			
2	8200	1	132			
1	11	0	2	0	
2	8201	1	132			
2	8202	1	137			
1	14	0	2	0	
2	8203	1	137			
2	8204	1	137			
1	17	0	2	0	
2	8205	1	137			
2	8206	1	137			
1	20	0	2	0	
2	8207	1	137			
2	8208	1	137			
1	23	0	1	0	
1	24	0	1	0	
1	25	0	1	0	
1	26	0	1	0	
1	27	0	3	0	
2	8211	1	137			
2	8212	1	137			
2	8222	1	141			
1	31	0	2	0	
2	8223	1	141			
2	8224	1	141			
1	34	0	2	0	
2	8227	1	146			
2	8228	1	146			
1	37	0	2	0	
2	8229	1	149			
2	8231	1	152			
1	40	0	2	0	
2	8232	1	152			
2	8233	1	155			
1	43	0	2	0	
2	8235	1	158			
2	8237	1	161			
1	46	0	2	0	
2	8239	1	164			
2	8240	1	164			
1	49	0	2	0	
2	8241	1	167			
2	8243	1	170			
1	52	0	1	0	
1	53	0	1	0	
1	54	0	7	0	
2	8245	1	173			
2	8244	1	170			
2	8246	1	173			
2	8242	1	167			
2	8249	1	179			
2	8250	1	179			
1	61	0	2	0	
2	8253	1	185			
2	8254	1	185			
1	64	0	2	0	
2	8257	1	191			
2	8251	1	182			
1	67	0	2	0	
2	8259	1	194			
2	8261	1	197			
1	70	0	2	0	
2	8263	1	200			
2	8255	1	188			
1	73	0	2	0	
2	8265	1	203			
2	8264	1	200			
1	76	0	2	0	
2	8266	1	203			
2	8262	1	197			
1	79	0	1	0	
1	80	0	1	0	
1	81	0	1	0	
1	82	0	1	0	
1	83	0	2	0	
2	8267	1	206			
2	8268	1	206			
1	86	0	1	0	
1	87	0	1	0	
1	88	0	2	0	
2	8278	1	210			
2	8279	1	210			
1	91	0	2	0	
2	8280	1	210			
2	8281	1	210			
1	94	0	2	0	
2	8282	1	210			
2	8283	1	210			
1	97	0	2	0	
2	8289	1	218			
2	8290	1	218			
1	100	0	2	0	
2	8291	1	218			
2	8292	1	218			
1	103	0	2	0	
2	8293	1	218			
2	8294	1	218			
1	106	0	2	0	
2	8295	1	218			
2	8300	1	226			
1	109	0	2	0	
2	8301	1	226			
2	8302	1	226			
2	8304	1	226			
1	112	0	1	0	
2	8306	1	226			
1	113	0	1	0	
1	114	0	1	0	
1	115	0	1	0	
1	116	0	1	0	
1	117	0	1	0	
1	118	0	1	0	
1	119	0	1	0	
1	120	0	1	0	
1	121	0	1	0	
1	122	0	1	0	
1	123	0	2	0	
2	8311	1	234			
2	8312	1	234			
1	126	0	1	0	
1	127	0	1	0	
1	128	0	1	0	
1	129	0	1	0	
1	130	0	1	0	
1	131	0	1	0	
1	132	0	2	0	
2	8322	1	242			
2	8323	1	242			
1	135	0	1	0	
1	136	0	1	0	
3	137	0	0	0	
2	8324	1	242			
2	8325	1	242			
1	140	0	1	0	
3	141	0	0	0	
2	8327	1	242			
2	8328	1	242			
1	145	0	1	0	
1	146	0	2	0	
2	8331	1	242			
1	149	0	2	0	
2	8342	1	245			
2	8334	1	242			
1	152	0	2	0	
2	8344	1	248			
2	8345	1	248			
1	155	0	2	0	
2	8346	1	248			
2	8347	1	248			
1	158	0	2	0	
2	8348	1	248			
2	8349	1	248			
1	161	0	2	0	
2	8350	1	248			
2	8351	1	248			
1	164	0	2	0	
2	8352	1	248			
2	8353	1	248			
1	167	0	2	0	
2	8354	1	248			
2	8355	1	248			
1	170	0	2	0	
2	8356	1	248			
2	8357	1	248			
1	173	0	2	0	
2	8358	1	248			
2	8361	1	248			
1	176	0	2	0	
2	8366	1	251			
2	8369	1	251			
1	179	0	2	0	
2	8370	1	251			
2	8372	1	251			
1	182	0	2	0	
2	8373	1	251			
2	8375	1	251			
1	185	0	2	0	
2	8376	1	251			
2	8371	1	251			
1	188	0	2	0	
2	8374	1	251			
2	8377	1	251			
1	191	0	2	0	
2	8378	1	251			
2	8379	1	251			
1	194	0	2	0	
2	8387	1	254			
2	8388	1	254			
1	197	0	2	0	
2	8389	1	254			
2	8390	1	254			
1	200	0	2	0	
2	8391	1	254			
2	8392	1	254			
1	203	0	2	0	
2	8393	1	254			
2	8394	1	254			
1	206	0	11	0	
2	8395	1	254			
2	8396	1	254			
1	209	0	1	0	
1	210	0	11	0	
2	8397	1	254			
2	8398	1	254			
2	8399	1	254			
2	8406	1	257			
2	8407	1	257			
2	8408	1	257			
1	217	0	1	0	
1	218	0	11	0	
2	8409	1	257			
2	8410	1	257			
2	8411	1	257			
2	8412	1	257			
2	8413	1	257			
2	8414	1	257			
1	225	0	1	0	
1	226	0	11	0	
2	8417	1	265			
2	8418	1	265			
2	8419	1	265			
2	8420	1	265			
2	8421	1	265			
2	8422	1	265			
1	233	0	1	0	
1	234	0	11	0	
2	8423	1	265			
2	8428	1	273			
2	8429	1	273			
2	8430	1	273			
2	8431	1	273			
2	8432	1	273			
1	241	0	1	0	
1	242	0	20	0	
2	8433	1	273			
2	8434	1	273			
1	245	0	2	0	
2	8435	1	273			
2	8439	1	281			
1	248	0	22	0	
2	8440	1	281			
2	8441	1	281			
1	251	0	21	0	
2	8442	1	281			
2	8443	1	281			
1	254	0	19	0	
2	8444	1	281			
2	8445	1	281			
1	257	0	11	0	
2	8446	1	281			
2	8447	1	281			
2	8450	1	289			
2	8453	1	293			
2	8454	1	293			
2	8455	1	293			
1	264	0	1	0	
1	265	0	11	0	
2	8456	1	293			
2	8457	1	293			
2	8460	1	299			
2	8458	1	293			
2	8462	1	302			
2	8463	1	302			
1	272	0	1	0	
1	273	0	11	0	
2	8464	1	302			
2	8465	1	302			
2	8466	1	302			
2	8469	1	308			
2	8470	1	308			
2	8471	1	308			
1	280	0	1	0	
1	281	0	11	0	
2	8472	1	308			
2	8473	1	308			
2	8474	1	308			
2	8475	1	308			
2	8476	1	308			
2	8477	1	308			
1	288	0	1	0	
1	289	0	3	0	
2	8480	1	316			
2	8481	1	316			
1	292	0	1	0	
3	293	0	0	0	
2	8482	1	316			
2	8483	1	316			
2	8484	1	316			
2	8485	1	316			
2	8486	1	316			
3	299	0	0	0	
2	8491	1	324			
2	8492	1	324			
1	302	0	7	0	
2	8493	1	324			
2	8494	1	324			
2	8495	1	324			
2	8496	1	324			
1	307	0	1	0	
1	308	0	11	0	
2	8501	1	332			
2	8502	1	332			
2	8503	1	332			
2	8504	1	332			
2	8505	1	332			
2	8506	1	332			
1	315	0	1	0	
1	316	0	11	0	
2	8507	1	332			
2	8508	1	332			
2	8509	1	332			
2	8510	1	332			
2	8513	1	335			
2	8514	1	335			
1	323	0	1	0	
1	324	0	10	0	
2	8515	1	335			
2	8516	1	335			
2	8517	1	335			
2	8518	1	335			
2	8519	1	335			
2	8520	1	335			
1	331	0	1	0	
1	332	0	12	0	
2	8525	1	338			
2	8521	1	335			
1	335	0	12	0	
2	8522	1	335			
2	8523	1	335			
1	338	0	2	0	
2	8524	1	335			
2	8527	1	341			
1	341	0	11	0	
2	8528	1	341			
2	8526	1	338			
2	8529	1	341			
2	8530	1	341			
2	8538	1	348			
2	8539	1	348			
1	348	0	2	0	
2	8540	1	351			
2	8541	1	351			
1	351	0	11	0	
2	8542	1	351			
2	8543	1	351			
2	8544	1	351			
2	8546	1	351			
2	8548	1	351			
2	8549	1	351			
1	358	0	2	0	
2	8551	1	358			
2	8552	1	358			
1	361	0	7	0	
2	8554	1	361			
2	8555	1	361			
2	8556	1	361			
2	8553	1	361			
1	366	0	2	0	
2	8557	1	361			
2	8560	1	366			
1	369	0	3	0	
2	8562	1	369			
2	8563	1	369			
2	8561	1	366			
1	372	0	1	0	
1	373	0	1	0	
1	374	0	13	0	
2	8565	1	374			
2	8566	1	374			
2	8567	1	374			
2	8568	1	374			
2	8569	1	374			
2	8570	1	374			
2	8571	1	374			
2	8572	1	374			
2	8573	1	374			
2	8574	1	374			
1	386	0	2	0	
2	8578	1	386			
2	8579	1	386			
1	389	0	12	0	
2	8580	1	389			
2	8581	1	389			
2	8582	1	389			
2	8583	1	389			
2	8584	1	389			
2	8585	1	389			
2	8586	1	389			
2	8587	1	389			
2	8588	1	389			
2	8589	1	389			
1	400	0	12	0	
2	8592	1	400			
2	8593	1	400			
2	8594	1	400			
2	8595	1	400			
2	8596	1	400			
2	8597	1	400			
2	8598	1	400			
2	8599	1	400			
2	8600	1	400			
2	8601	1	400			
1	411	0	12	0	
2	8604	1	411			
2	8605	1	411			
2	8606	1	411			
2	8607	1	411			
2	8608	1	411			
2	8609	1	411			
2	8610	1	411			
2	8611	1	411			
2	8612	1	411			
2	8613	1	411			
1	422	0	14	0	
2	8225	1	141			
2	8616	1	422			
2	8617	1	422			
2	8618	1	422			
2	8619	1	422			
2	8620	1	422			
2	8621	1	422			
2	8622	1	422			
2	8623	1	422			
2	8624	1	422			
2	8625	1	422			
2	8626	1	422			
1	435	0	12	0	
2	8627	1	422			
2	8226	1	141			
2	8630	1	435			
2	8631	1	435			
2	8632	1	435			
2	8633	1	435			
2	8634	1	435			
2	8635	1	435			
2	8636	1	435			
2	8637	1	435			
1	446	0	12	0	
2	8638	1	435			
2	8230	1	149			
2	8639	1	435			
2	8642	1	446			
2	8643	1	446			
2	8644	1	446			
2	8645	1	446			
2	8646	1	446			
2	8647	1	446			
2	8648	1	446			
1	457	0	12	0	
2	8649	1	446			
2	8650	1	446			
2	8651	1	446			
2	8652	1	446			
2	8654	1	457			
2	8655	1	457			
2	8656	1	457			
2	8657	1	457			
2	8658	1	457			
2	8659	1	457			
1	468	0	12	0	
2	8234	1	155			
2	8660	1	457			
2	8661	1	457			
2	8662	1	457			
2	8663	1	457			
2	8666	1	468			
2	8667	1	468			
2	8668	1	468			
2	8669	1	468			
2	8236	1	158			
1	479	0	12	0	
2	8670	1	468			
2	8671	1	468			
2	8672	1	468			
2	8673	1	468			
2	8674	1	468			
2	8675	1	468			
2	8678	1	479			
2	8679	1	479			
2	8238	1	161			
2	8680	1	479			
1	490	0	14	0	
2	8681	1	479			
2	8682	1	479			
2	8683	1	479			
2	8684	1	479			
2	8685	1	479			
2	8686	1	479			
2	8687	1	479			
2	8690	1	490			
2	8691	1	490			
2	8692	1	490			
2	8693	1	490			
2	8694	1	490			
1	503	0	12	0	
2	8695	1	490			
2	8696	1	490			
2	8697	1	490			
2	8698	1	490			
2	8699	1	490			
2	8700	1	490			
2	8701	1	490			
2	8702	1	490			
2	8704	1	503			
2	8705	1	503			
1	514	0	10	0	
2	8706	1	503			
2	8707	1	503			
2	8708	1	503			
2	8709	1	503			
2	8710	1	503			
2	8711	1	503			
2	8712	1	503			
2	8713	1	503			
1	523	0	12	0	
2	8716	1	514			
2	8717	1	514			
2	8718	1	514			
2	8719	1	514			
2	8720	1	514			
2	8721	1	514			
2	8722	1	514			
2	8723	1	514			
2	8724	1	514			
2	8247	1	176			
1	534	0	12	0	
2	8726	1	523			
2	8727	1	523			
2	8728	1	523			
2	8730	1	523			
2	8731	1	523			
2	8729	1	523			
2	8248	1	176			
2	8732	1	523			
2	8733	1	523			
2	8734	1	523			
1	545	0	3	0	
2	8738	1	534			
2	8739	1	534			
2	8740	1	534			
3	549	0	0	0	
2	8741	1	534			
2	8742	1	534			
1	552	0	3	0	
2	8743	1	534			
2	8744	1	534			
2	8745	1	534			
1	556	0	2	0	
2	8746	1	534			
2	8750	1	545			
1	559	0	2	0	
2	8752	1	545			
2	8753	1	549			
1	562	0	3	0	
2	8755	1	552			
2	8751	1	545			
2	8756	1	552			
1	566	0	4	0	
2	8758	1	556			
2	8760	1	559			
2	8761	1	559			
2	8762	1	562			
1	571	0	22	0	
2	8763	1	562			
2	8759	1	556			
1	574	0	22	0	
2	8765	1	566			
2	8764	1	562			
1	577	0	22	0	
2	8769	1	571			
2	8770	1	571			
1	580	0	22	0	
2	8771	1	571			
2	8772	1	571			
1	583	0	4	0	
2	8773	1	571			
2	8774	1	571			
2	8775	1	571			
2	8776	1	571			
1	588	0	10	0	
2	8777	1	571			
2	8778	1	571			
1	591	0	1	0	
3	592	0	0	0	
2	8779	1	571			
2	8780	1	571			
1	595	0	1	0	
1	596	0	1	0	
1	597	0	1	0	
1	598	0	1	0	
1	599	0	3	0	
2	8791	1	574			
2	8792	1	574			
2	8793	1	574			
1	603	0	3	0	
2	8794	1	574			
2	8795	1	574			
2	8796	1	574			
1	607	0	22	0	
2	8797	1	574			
2	8798	1	574			
1	610	0	22	0	
2	8799	1	574			
2	8800	1	574			
1	613	0	22	0	
2	8801	1	574			
2	8802	1	574			
1	616	0	22	0	
2	8803	1	574			
2	8804	1	574			
1	619	0	29	0	
2	8805	1	574			
2	8813	1	577			
2	8814	1	577			
2	8815	1	577			
2	8816	1	577			
1	625	0	31	0	
2	8817	1	577			
2	8818	1	577			
2	8819	1	577			
2	8820	1	577			
2	8821	1	577			
1	631	0	1	0	
2	8822	1	577			
2	8823	1	577			
2	8824	1	577			
2	8825	1	577			
2	8826	1	577			
2	8827	1	577			
2	8828	1	577			
2	8829	1	577			
2	8830	1	577			
2	8831	1	577			
2	8832	1	577			
2	8835	1	580			
2	8836	1	580			
2	8837	1	580			
2	8838	1	580			
2	8839	1	580			
2	8840	1	580			
2	8841	1	580			
2	8842	1	580			
2	8843	1	580			
2	8844	1	580			
2	8845	1	580			
2	8846	1	580			
2	8847	1	580			
2	8848	1	580			
2	8849	1	580			
2	8850	1	580			
2	8851	1	580			
2	8852	1	580			
2	8853	1	580			
2	8854	1	580			
2	8855	1	580			
2	8856	1	580			
2	8857	1	583			
2	8272	1	206			
2	8273	1	206			
2	9902	1	5389			
2	8861	1	588			
2	8862	1	588			
2	8863	1	588			
2	8864	1	588			
2	8865	1	588			
2	8866	1	588			
2	8274	1	206			
2	8275	1	206			
2	8867	1	588			
2	8868	1	588			
2	8871	1	599			
2	8872	1	599			
2	8276	1	206			
2	8874	1	603			
2	8869	1	588			
2	8277	1	206			
2	8877	1	607			
2	8878	1	607			
2	8879	1	607			
2	8880	1	607			
2	8881	1	607			
2	8882	1	607			
2	8883	1	607			
2	8884	1	607			
2	8885	1	607			
2	8886	1	607			
2	8887	1	607			
2	8888	1	607			
2	8889	1	607			
2	8890	1	607			
2	8891	1	607			
2	8892	1	607			
2	8893	1	607			
2	8894	1	607			
2	8895	1	607			
2	8896	1	607			
2	8897	1	607			
2	8898	1	607			
2	8899	1	610			
2	8900	1	610			
2	8901	1	610			
2	8902	1	610			
2	8903	1	610			
2	8904	1	610			
2	8905	1	610			
2	8906	1	610			
2	8907	1	610			
2	8908	1	610			
2	8909	1	610			
2	8910	1	610			
2	8284	1	210			
2	8911	1	610			
2	8912	1	610			
2	8913	1	610			
2	8914	1	610			
2	8285	1	210			
2	8915	1	610			
2	8916	1	610			
2	8917	1	610			
2	8918	1	610			
2	8921	1	613			
2	8922	1	613			
2	8923	1	613			
2	8924	1	613			
2	8925	1	613			
2	8926	1	613			
2	8927	1	613			
2	8928	1	613			
2	8929	1	613			
2	8930	1	613			
2	8931	1	613			
2	8932	1	613			
2	8287	1	210			
2	8288	1	210			
2	8933	1	613			
2	8934	1	613			
2	8935	1	613			
2	8936	1	613			
2	8937	1	613			
2	8938	1	613			
2	8939	1	613			
2	8940	1	613			
2	8943	1	616			
2	8944	1	616			
2	8945	1	616			
2	8946	1	616			
2	8947	1	616			
2	8948	1	616			
2	8949	1	616			
2	8950	1	616			
2	8951	1	616			
2	8952	1	616			
2	8953	1	616			
2	8954	1	616			
2	8955	1	616			
2	8956	1	616			
2	8957	1	616			
2	8958	1	616			
2	8959	1	616			
2	8960	1	616			
2	8961	1	616			
2	8962	1	616			
2	8963	1	616			
2	8964	1	616			
2	8965	1	619			
2	8966	1	619			
2	8967	1	619			
2	8968	1	619			
2	8969	1	619			
2	8970	1	619			
2	8971	1	619			
2	8296	1	218			
2	8972	1	619			
2	8973	1	619			
2	8974	1	619			
2	8975	1	619			
2	8297	1	218			
2	8976	1	619			
2	8977	1	619			
2	8978	1	619			
2	8979	1	619			
2	8298	1	218			
2	8980	1	619			
2	8981	1	619			
2	8982	1	619			
2	8983	1	619			
2	8299	1	218			
2	8984	1	619			
2	8985	1	619			
2	8986	1	619			
2	8987	1	619			
2	8988	1	619			
2	8989	1	619			
2	8994	1	625			
2	8995	1	625			
2	8996	1	625			
2	8997	1	625			
2	8998	1	625			
2	8999	1	625			
2	9000	1	625			
2	9001	1	625			
2	9002	1	625			
2	9003	1	625			
2	9004	1	625			
2	9005	1	625			
2	9006	1	625			
2	8303	1	226			
2	9007	1	625			
2	9008	1	625			
2	9009	1	625			
2	9010	1	625			
2	9011	1	625			
2	9012	1	625			
2	9013	1	625			
2	9014	1	625			
2	9015	1	625			
2	8305	1	226			
2	9016	1	625			
2	9017	1	625			
2	9018	1	625			
2	9019	1	625			
2	9020	1	625			
2	9021	1	625			
2	9022	1	625			
2	9025	1	1067			
2	9026	1	1067			
2	8307	1	226			
2	9027	1	1067			
2	9028	1	1067			
2	9029	1	1067			
2	9030	1	1067			
2	9031	1	1067			
2	9032	1	1067			
2	9033	1	1067			
2	9034	1	1067			
2	9035	1	1067			
2	9036	1	1067			
2	9037	1	1080			
2	9038	1	1080			
2	9040	1	1080			
2	9041	1	1080			
2	9042	1	1080			
2	9043	1	1080			
2	9044	1	1080			
2	9045	1	1080			
2	9046	1	1080			
2	9047	1	1080			
2	9048	1	1092			
2	9049	1	1092			
2	9050	1	1092			
2	9051	1	1092			
2	9052	1	1092			
2	9053	1	1092			
2	9054	1	1092			
2	9055	1	1092			
2	9056	1	1092			
2	9057	1	1092			
2	9058	1	1092			
2	8313	1	234			
2	9059	1	1104			
2	9060	1	1104			
2	9061	1	1104			
2	9062	1	1104			
2	9063	1	1104			
2	8314	1	234			
2	9064	1	1104			
2	9065	1	1104			
2	9066	1	1104			
2	9067	1	1104			
2	9068	1	1104			
2	9069	1	1104			
2	9070	1	1104			
2	8315	1	234			
2	8316	1	234			
2	9071	1	1157			
2	9072	1	1157			
2	9077	1	1475			
2	9078	1	1475			
2	9079	1	1475			
2	8317	1	234			
2	9080	1	1583			
2	8318	1	234			
2	9081	1	1583			
2	9084	1	1588			
2	9085	1	1588			
2	9086	1	1588			
2	8319	1	234			
2	9088	1	1588			
2	9087	1	1588			
2	9089	1	1660			
2	9090	1	1660			
2	9083	1	1583			
2	8320	1	234			
2	9091	1	1660			
2	9095	1	1758			
2	9096	1	1758			
2	9097	1	2653			
2	9098	1	2653			
2	9099	1	2653			
2	9100	1	2653			
2	9101	1	2653			
2	8321	1	234			
2	9094	1	1755			
2	9102	1	2653			
2	9103	1	2653			
2	9104	1	2653			
2	9107	1	2664			
2	9108	1	2664			
2	9109	1	2664			
2	9110	1	2664			
2	9111	1	2664			
2	9112	1	2664			
2	9105	1	2653			
2	9113	1	2664			
2	9114	1	2664			
2	9115	1	2664			
2	9117	1	2681			
2	9118	1	2681			
2	9119	1	2681			
2	9120	1	2681			
2	9121	1	2681			
2	9122	1	2681			
2	8326	1	242			
2	9123	1	2681			
2	9124	1	2681			
2	9125	1	2681			
2	9127	1	2692			
2	9128	1	2692			
2	9129	1	2692			
2	9130	1	2692			
2	9131	1	2692			
2	9132	1	2692			
2	9133	1	2692			
2	9134	1	2692			
2	9155	1	2739			
2	9135	1	2692			
2	9137	1	2728			
2	8329	1	242			
2	9138	1	2728			
2	9139	1	2728			
2	9140	1	2728			
2	9141	1	2728			
2	8330	1	242			
2	9142	1	2728			
2	9143	1	2728			
2	9144	1	2728			
2	9959	1	5441			
2	9147	1	2739			
2	9148	1	2739			
2	9149	1	2739			
2	9150	1	2739			
2	9151	1	2739			
2	8332	1	242			
2	9152	1	2739			
2	9153	1	2739			
2	9154	1	2739			
2	9157	1	2756			
2	8333	1	242			
2	9158	1	2756			
2	9159	1	2756			
2	9160	1	2756			
2	9161	1	2756			
2	9162	1	2756			
2	9163	1	2756			
2	9164	1	2756			
2	9165	1	2756			
2	9167	1	2767			
2	8335	1	242			
2	9168	1	2767			
2	9169	1	2767			
2	9170	1	2767			
2	9171	1	2767			
2	8336	1	242			
2	9172	1	2767			
2	9173	1	2767			
2	9174	1	2767			
2	9177	1	2779			
2	8337	1	242			
2	9178	1	2779			
2	9179	1	2779			
2	9180	1	2779			
2	9181	1	2779			
2	8338	1	242			
2	9182	1	2779			
2	9183	1	2779			
2	9184	1	2779			
2	9187	1	2790			
2	8339	1	242			
2	9188	1	2790			
2	9189	1	2790			
2	9190	1	2790			
2	9191	1	2790			
2	8340	1	242			
2	9185	1	2779			
2	9192	1	2790			
2	9193	1	2790			
2	9197	1	2801			
2	9198	1	2801			
2	9199	1	2801			
2	9200	1	2801			
2	9201	1	2801			
2	8341	1	242			
2	9202	1	2801			
2	9203	1	2801			
2	9204	1	2801			
2	9205	1	2801			
2	9207	1	2812			
2	9208	1	2812			
2	9209	1	2812			
2	9210	1	2812			
2	9211	1	2812			
2	9212	1	2812			
2	9213	1	2812			
2	9214	1	2812			
2	8343	1	245			
2	9215	1	2812			
2	9217	1	2855			
2	9218	1	2855			
2	9219	1	2855			
2	9220	1	2855			
2	9221	1	2855			
2	9222	1	2861			
2	9223	1	2861			
2	9224	1	2861			
2	9225	1	2861			
2	9226	1	2861			
2	9227	1	2882			
2	9228	1	2882			
2	9229	1	2882			
2	9230	1	2882			
2	9231	1	2882			
2	9232	1	2882			
2	9233	1	2882			
0	1042	7	1	2	135	631	
0	1043	5	1	1	591	
2	9235	1	2891			
2	9236	1	2891			
2	9237	1	2891			
2	9238	1	2891			
2	9239	1	2891			
2	9240	1	2891			
2	9241	1	2891			
2	9242	1	2891			
2	9243	1	2891			
2	9244	1	2942			
2	9245	1	2942			
2	9246	1	2942			
2	9247	1	2942			
2	9249	1	2948			
2	9250	1	2948			
2	9251	1	2948			
2	9252	1	2948			
2	9253	1	2948			
2	9248	1	2942			
2	9254	1	2964			
2	9255	1	2964			
2	9256	1	2964			
2	9258	1	3041			
0	1067	5	12	1	595	
2	9259	1	3041			
2	9260	1	3041			
2	9261	1	3041			
2	9262	1	3041			
2	9257	1	2964			
2	9263	1	3041			
2	9264	1	3041			
2	9265	1	3041			
2	9268	1	3052			
2	9269	1	3052			
2	9270	1	3052			
2	9271	1	3052			
0	1080	5	11	1	596	
2	9272	1	3052			
2	9273	1	3052			
2	9266	1	3041			
2	9274	1	3052			
2	9275	1	3052			
2	9276	1	3052			
2	9277	1	3052			
2	9984	1	5470			
2	9278	1	3063			
2	9282	1	3068			
2	9283	1	3068			
0	1092	5	11	1	597	
2	9284	1	3075			
2	9285	1	3075			
2	9286	1	3075			
2	9287	1	3075			
2	8359	1	248			
2	9288	1	3075			
2	9289	1	3075			
2	9290	1	3075			
2	9291	1	3075			
2	8360	1	248			
2	9294	1	3086			
0	1104	5	12	1	598	
2	9295	1	3086			
2	9296	1	3086			
2	9297	1	3086			
2	9298	1	3086			
2	9299	1	3086			
2	9300	1	3086			
2	9301	1	3086			
2	8362	1	248			
2	9304	1	3097			
2	9305	1	3097			
2	9306	1	3097			
2	9307	1	3097			
2	8363	1	248			
2	9308	1	3097			
2	9309	1	3097			
2	9310	1	3097			
2	9311	1	3097			
2	8364	1	248			
2	9314	1	3108			
2	9315	1	3108			
2	9316	1	3108			
2	9312	1	3097			
2	8365	1	248			
2	9317	1	3108			
2	9318	1	3108			
2	9319	1	3108			
2	9320	1	3108			
2	9324	1	3119			
2	9325	1	3119			
2	9326	1	3119			
2	9327	1	3119			
2	9328	1	3119			
3	1137	5	0	1	8750	
3	1138	5	0	1	8538	
3	1139	5	0	1	8560	
3	1140	7	0	2	8755	8762	
3	1141	5	0	1	8753	
3	1142	5	0	1	8751	
3	1143	5	0	1	8752	
3	1144	5	0	1	8525	
3	1145	5	0	1	8551	
0	1146	6	1	2	373	1	
3	1147	7	0	2	8222	145	
0	1148	5	1	1	592	
0	1149	5	1	1	1042	
0	1150	7	1	2	1043	8144	
0	1151	7	1	2	8578	8758	
3	1152	5	0	1	8342	
3	1153	5	0	1	8756	
3	1154	5	0	1	8763	
3	1155	5	0	1	8760	
0	1156	7	1	4	8579	8761	8759	8757	
0	1157	5	3	1	8765	
2	9344	1	3147			
2	9345	1	3147			
2	9346	1	3147			
2	9347	1	3147			
2	9348	1	3147			
2	9349	1	3147			
2	9354	1	3158			
2	9350	1	3147			
2	9355	1	3158			
2	9351	1	3147			
2	9356	1	3158			
2	9352	1	3147			
2	9357	1	3158			
2	9358	1	3158			
2	9364	1	3169			
2	9365	1	3169			
2	9366	1	3169			
2	9367	1	3169			
2	9368	1	3169			
2	9369	1	3169			
2	9370	1	3169			
2	9371	1	3169			
2	9372	1	3169			
2	9373	1	3169			
2	9374	1	3180			
2	9375	1	3180			
2	9376	1	3180			
2	9377	1	3180			
2	9378	1	3180			
2	9379	1	3180			
2	9380	1	3180			
2	9381	1	3180			
2	9382	1	3180			
2	9383	1	3180			
2	9384	1	3456			
2	9385	1	3456			
2	9386	1	3691			
2	9387	1	3691			
2	9388	1	3691			
2	9389	1	3691			
2	9390	1	3691			
2	9391	1	3691			
2	9392	1	3691			
2	9393	1	3691			
2	8380	1	251			
2	9394	1	3705			
2	9395	1	3705			
2	9397	1	3732			
2	9398	1	3732			
2	8381	1	251			
2	9399	1	3732			
2	9400	1	3732			
2	9401	1	3732			
2	9402	1	3732			
2	8382	1	251			
2	9405	1	3771			
2	9406	1	3771			
2	9403	1	3732			
2	9408	1	3775			
2	8383	1	251			
2	9409	1	3775			
0	1219	5	3	1	8857	
2	9411	1	3789			
2	9410	1	3775			
2	9414	1	3793			
2	8384	1	251			
2	9407	1	3771			
2	9417	1	3797			
2	9418	1	3797			
2	9415	1	3793			
2	8385	1	251			
2	9421	1	3810			
2	9422	1	3810			
2	9423	1	3813			
2	9424	1	3813			
2	8386	1	251			
2	9425	1	3816			
2	9427	1	3819			
2	9419	1	3797			
2	9429	1	3824			
2	9428	1	3819			
2	9431	1	3842			
2	9432	1	3842			
2	9433	1	3842			
2	9434	1	3842			
2	9435	1	3842			
2	9436	1	3842			
2	9437	1	3842			
2	9438	1	3842			
2	9430	1	3824			
2	9440	1	3849			
2	9441	1	3849			
2	9442	1	3849			
2	9443	1	3849			
2	9444	1	3849			
2	9445	1	3849			
2	9446	1	3849			
2	9439	1	3842			
2	9448	1	3855			
2	9449	1	3855			
2	9450	1	3855			
2	9451	1	3855			
2	9452	1	3855			
2	9453	1	3855			
2	9454	1	3855			
2	9447	1	3849			
2	9456	1	3861			
2	9457	1	3861			
2	9458	1	3861			
2	9459	1	3861			
2	9460	1	3861			
2	9461	1	3861			
2	9462	1	3861			
2	9455	1	3855			
2	9464	1	3867			
2	9465	1	3867			
2	9466	1	3867			
2	9467	1	3867			
2	9468	1	3867			
2	9469	1	3867			
2	9470	1	3867			
2	9471	1	3867			
2	9472	1	3873			
2	9473	1	3873			
2	9474	1	3873			
2	9475	1	3873			
2	9476	1	3873			
2	9477	1	3873			
2	9478	1	3873			
2	9479	1	3873			
2	9480	1	3873			
2	9481	1	3873			
2	9482	1	3881			
2	9483	1	3881			
2	9484	1	3881			
2	9485	1	3881			
2	9486	1	3881			
2	9487	1	3881			
2	9488	1	3881			
2	9489	1	3881			
2	9490	1	3887			
2	9491	1	3887			
2	9492	1	3887			
2	9493	1	3887			
2	9494	1	3887			
2	8400	1	254			
2	9495	1	3887			
2	9496	1	3887			
2	9498	1	3893			
2	9499	1	3893			
2	8401	1	254			
2	9500	1	3893			
2	9501	1	3893			
2	9502	1	3893			
2	9503	1	3893			
2	8402	1	254			
2	9506	1	3911			
2	9507	1	3911			
2	9508	1	3921			
2	9509	1	3921			
2	8403	1	254			
2	9510	1	3921			
2	9511	1	3921			
2	9504	1	3893			
2	9505	1	3893			
2	8404	1	254			
2	9512	1	3921			
2	9513	1	3921			
2	9514	1	3921			
2	9515	1	3921			
2	8405	1	254			
2	9516	1	3921			
2	9517	1	3921			
2	9518	1	3921			
2	9519	1	3921			
2	9525	1	3927			
2	9526	1	3927			
2	9527	1	3927			
2	9528	1	3927			
2	9529	1	3927			
2	9530	1	3927			
2	9531	1	3927			
2	9532	1	3927			
2	9533	1	3933			
2	9534	1	3933			
2	9535	1	3933			
2	9536	1	3933			
2	9537	1	3933			
2	9538	1	3933			
2	9539	1	3933			
2	9540	1	3933			
2	9541	1	3942			
2	9542	1	3942			
2	9543	1	3942			
2	9544	1	3942			
2	9545	1	3942			
2	9546	1	3942			
2	9547	1	3942			
2	9548	1	3942			
2	9549	1	3948			
2	9550	1	3948			
2	9551	1	3948			
2	9552	1	3948			
2	9553	1	3948			
2	9554	1	3948			
2	9555	1	3948			
2	9556	1	3948			
2	9557	1	3948			
2	9558	1	3948			
2	9559	1	3956			
2	9560	1	3956			
2	9561	1	3956			
2	9562	1	3956			
2	9563	1	3956			
2	9564	1	3956			
2	9565	1	3956			
2	9566	1	3956			
2	9567	1	3962			
2	9568	1	3962			
2	9569	1	3962			
2	8415	1	257			
2	9570	1	3962			
2	9571	1	3962			
2	9572	1	3962			
2	9573	1	3962			
2	9574	1	3962			
2	8416	1	257			
2	9577	1	3968			
2	9578	1	3968			
2	9579	1	3968			
2	9580	1	3968			
2	9581	1	3968			
2	9582	1	3968			
2	9583	1	3968			
2	9584	1	3968			
2	9585	1	3984			
2	9586	1	3984			
2	9587	1	4008			
2	9588	1	4008			
2	9589	1	4011			
2	9590	1	4011			
2	9591	1	4021			
2	9592	1	4021			
2	9593	1	4067			
2	9594	1	4067			
2	9595	1	4080			
2	9596	1	4080			
2	9597	1	4080			
2	9598	1	4088			
2	9599	1	4088			
2	9600	1	4091			
2	9601	1	4091			
2	9602	1	4094			
2	9603	1	4094			
2	9604	1	4097			
2	9605	1	4097			
2	9606	1	4100			
2	9607	1	4100			
2	9608	1	4103			
2	9609	1	4103			
2	9610	1	4106			
2	9611	1	4106			
2	9612	1	4109			
2	9613	1	4109			
2	9614	1	4144			
2	9615	1	4144			
2	8424	1	265			
2	9616	1	4147			
2	9618	1	4153			
2	9619	1	4153			
2	9620	1	4156			
2	8425	1	265			
2	9622	1	4159			
2	9623	1	4159			
2	9624	1	4188			
2	9625	1	4188			
2	8426	1	265			
2	9626	1	4191			
2	9627	1	4191			
2	9621	1	4156			
2	9630	1	4203			
2	8427	1	265			
2	9632	1	4225			
2	9628	1	4200			
2	9634	1	4228			
2	9635	1	4228			
2	9636	1	4231			
2	9633	1	4225			
2	9638	1	4234			
2	9639	1	4234			
2	9640	1	4237			
2	9637	1	4231			
2	9642	1	4240			
2	9643	1	4240			
2	9644	1	4243			
2	9641	1	4237			
2	9646	1	4246			
2	9647	1	4246			
2	9648	1	4249			
2	9649	1	4249			
2	9650	1	4252			
2	9651	1	4252			
2	9652	1	4255			
2	9653	1	4255			
2	9654	1	4258			
2	9655	1	4258			
2	9656	1	4264			
2	9657	1	4264			
2	9658	1	4280			
2	9659	1	4280			
2	9660	1	4280			
2	9661	1	4284			
2	9662	1	4284			
2	9663	1	4284			
2	9664	1	4284			
2	9665	1	4284			
2	9666	1	4290			
0	1475	7	3	2	8145	8147	
2	9667	1	4290			
2	9668	1	4290			
2	9669	1	4290			
2	9670	1	4290			
2	9671	1	4290			
2	9673	1	4298			
2	9674	1	4298			
2	9675	1	4301			
2	8436	1	273			
2	9676	1	4301			
2	9678	1	4305			
2	9679	1	4305			
2	9680	1	4305			
2	8437	1	273			
2	9682	1	4310			
2	9683	1	4310			
2	9684	1	4310			
2	9685	1	4310			
2	8438	1	273			
2	9687	1	4316			
2	9681	1	4305			
2	9686	1	4310			
2	9690	1	4320			
2	9691	1	4320			
2	9692	1	4320			
2	9693	1	4320			
2	9694	1	4325			
2	9695	1	4325			
2	9696	1	4325			
2	9697	1	4325			
2	9698	1	4325			
2	9699	1	4325			
2	9700	1	4332			
2	9701	1	4332			
2	9702	1	4332			
2	9703	1	4336			
2	9704	1	4336			
2	9705	1	4336			
2	9706	1	4336			
2	9707	1	4336			
2	9708	1	4342			
2	9709	1	4342			
2	9710	1	4342			
2	9711	1	4342			
2	9712	1	4342			
2	9713	1	4342			
2	9714	1	4349			
2	9715	1	4349			
2	9716	1	4349			
2	9717	1	4349			
2	9718	1	4349			
2	9719	1	4349			
2	9720	1	4349			
2	9721	1	4349			
2	9722	1	4357			
2	9723	1	4357			
2	9724	1	4357			
2	9725	1	4357			
2	9726	1	4357			
2	9727	1	4357			
2	9728	1	4357			
2	9729	1	4357			
2	9730	1	4364			
2	9731	1	4364			
2	9732	1	4364			
2	9733	1	4364			
2	9734	1	4364			
2	9735	1	4364			
2	9736	1	4364			
2	8448	1	281			
2	9737	1	4364			
2	9738	1	4364			
2	9739	1	4364			
2	9740	1	4364			
2	8449	1	281			
2	9742	1	4379			
2	9743	1	4379			
2	9744	1	4379			
2	9745	1	4379			
2	9747	1	4385			
2	9748	1	4385			
2	9749	1	4385			
2	9750	1	4385			
2	9751	1	4385			
2	8451	1	289			
2	9752	1	4385			
2	9754	1	4396			
2	9755	1	4396			
2	9756	1	4396			
2	8452	1	289			
2	9757	1	4400			
2	9758	1	4400			
2	9759	1	4400			
2	9761	1	4405			
2	9762	1	4405			
2	9763	1	4405			
2	9764	1	4405			
2	9765	1	4405			
2	9766	1	4405			
2	9767	1	4405			
2	9768	1	4418			
2	9769	1	4418			
2	9770	1	4418			
2	9771	1	4418			
2	9772	1	4418			
2	9773	1	4418			
2	10157	1	5655			
0	1583	7	4	2	8148	8146	
2	9776	1	4425			
2	9777	1	4425			
2	9778	1	4425			
2	9779	1	4425			
0	1588	5	5	1	8861	
2	9780	1	4425			
2	9781	1	4425			
2	9782	1	4425			
2	9783	1	4425			
2	9784	1	4425			
2	9785	1	4425			
2	9832	1	4646			
2	9788	1	4440			
2	9789	1	4440			
2	9790	1	4440			
2	9791	1	4440			
2	8459	1	293			
2	9792	1	4445			
2	9793	1	4445			
2	9794	1	4445			
2	9795	1	4445			
2	9796	1	4445			
2	9798	1	4456			
2	9799	1	4456			
2	9800	1	4456			
2	9801	1	4456			
2	8461	1	299			
2	9803	1	4462			
2	9804	1	4462			
2	9805	1	4462			
2	9806	1	4462			
2	9807	1	4462			
2	9808	1	4462			
2	9809	1	4477			
2	9810	1	4477			
2	9811	1	4477			
2	9812	1	4477			
2	9813	1	4477			
2	9814	1	4477			
2	9815	1	4477			
2	9816	1	4477			
2	9817	1	4524			
2	9818	1	4524			
2	9819	1	4524			
2	9820	1	4532			
2	9821	1	4532			
2	9822	1	4532			
2	9823	1	4575			
2	9824	1	4575			
2	9825	1	4605			
2	9826	1	4605			
2	9827	1	4608			
2	9828	1	4608			
2	9829	1	4627			
2	9830	1	4627			
2	9831	1	4646			
2	8467	1	302			
2	9833	1	4939			
2	9834	1	4939			
2	9835	1	4939			
2	9836	1	5049			
2	8468	1	302			
2	9837	1	5049			
2	9838	1	5150			
2	9840	1	5157			
2	9839	1	5150			
2	9842	1	5166			
2	9843	1	5166			
2	9844	1	5236			
2	9845	1	5236			
2	9846	1	5264			
2	9847	1	5264			
2	9848	1	5264			
2	9849	1	5264			
2	9850	1	5264			
2	9851	1	5264			
0	1660	5	4	1	8491	
2	9852	1	5264			
2	9853	1	5264			
2	9854	1	5264			
2	9856	1	5284			
2	9857	1	5284			
2	9858	1	5284			
2	9859	1	5284			
2	9860	1	5284			
2	9861	1	5284			
2	9862	1	5284			
2	9863	1	5284			
2	9864	1	5284			
2	9865	1	5284			
2	9866	1	5284			
2	9867	1	5284			
2	9868	1	5284			
2	10173	1	5671			
2	9869	1	5284			
2	9871	1	5315			
2	9872	1	5315			
2	9873	1	5315			
2	9874	1	5319			
2	9875	1	5319			
2	9876	1	5319			
2	9877	1	5319			
2	9878	1	5324			
2	9879	1	5324			
2	9880	1	5324			
2	9881	1	5328			
2	9882	1	5328			
2	9883	1	5328			
2	9884	1	5328			
2	9885	1	5346			
2	9886	1	5346			
2	8478	1	308			
2	9887	1	5371			
2	9888	1	5371			
2	9889	1	5377			
2	9891	1	5382			
2	8479	1	308			
2	9893	1	5385			
2	9892	1	5382			
2	9895	1	5389			
2	9896	1	5389			
2	9897	1	5389			
2	9898	1	5389			
2	9894	1	5385			
2	9899	1	5389			
2	9900	1	5389			
2	9901	1	5389			
2	9903	1	5396			
2	9904	1	5396			
2	9905	1	5396			
2	9906	1	5396			
2	9907	1	5396			
2	9908	1	5396			
2	9909	1	5396			
2	9910	1	5396			
2	9911	1	5396			
2	9912	1	5396			
2	9913	1	5396			
2	9914	1	5396			
2	9915	1	5407			
2	9916	1	5407			
2	9917	1	5407			
2	9918	1	5407			
2	9919	1	5407			
2	9920	1	5407			
2	9921	1	5407			
2	9922	1	5407			
2	9923	1	5407			
2	9924	1	5407			
2	9925	1	5407			
2	9926	1	5407			
2	9927	1	5418			
2	9928	1	5418			
2	9929	1	5418			
2	9930	1	5418			
2	9931	1	5418			
2	9932	1	5424			
2	8487	1	316			
2	9933	1	5424			
2	9934	1	5424			
2	9935	1	5424			
2	9936	1	5424			
2	8488	1	316			
2	9939	1	5431			
2	9940	1	5431			
2	9941	1	5431			
2	9942	1	5431			
2	8489	1	316			
2	9943	1	5431			
2	9944	1	5431			
2	9945	1	5431			
0	1755	5	2	1	8871	
2	8490	1	316			
2	9949	1	5441			
0	1758	5	2	1	8874	
2	9950	1	5441			
2	9951	1	5441			
2	9952	1	5441			
2	9953	1	5441			
2	9954	1	5441			
2	9955	1	5441			
2	9956	1	5441			
2	9957	1	5441			
2	9958	1	5441			
2	9960	1	5452			
2	9961	1	5452			
2	9962	1	5452			
2	9963	1	5452			
2	9964	1	5452			
2	9965	1	5452			
2	9966	1	5452			
2	9967	1	5452			
2	9968	1	5452			
2	9969	1	5452			
2	9970	1	5462			
2	9971	1	5462			
2	9972	1	5462			
2	9973	1	5462			
2	9974	1	5462			
2	9975	1	5462			
2	9976	1	5462			
2	9977	1	5470			
2	9978	1	5470			
2	9979	1	5470			
2	9980	1	5470			
2	9981	1	5470			
2	9982	1	5470			
2	8497	1	324			
2	9983	1	5470			
2	9985	1	5477			
2	9986	1	5477			
2	9987	1	5477			
2	8498	1	324			
2	9988	1	5477			
2	9989	1	5477			
2	9990	1	5477			
2	9991	1	5477			
2	8499	1	324			
2	9992	1	5477			
2	9993	1	5477			
2	9994	1	5477			
2	9997	1	5488			
2	8500	1	324			
2	9998	1	5488			
2	9999	1	5488			
2	10000	1	5488			
2	10001	1	5488			
2	10002	1	5488			
2	10003	1	5488			
2	10004	1	5488			
2	10005	1	5488			
2	9841	1	5157			
2	10008	1	5498			
2	10009	1	5498			
2	10010	1	5498			
2	10011	1	5498			
2	10012	1	5498			
2	10013	1	5498			
2	10014	1	5498			
2	8213	1	137			
2	10007	1	5488			
2	10017	1	5506			
2	10018	1	5506			
2	10019	1	5506			
2	10020	1	5506			
2	10021	1	5506			
2	10022	1	5506			
2	10023	1	5506			
2	10024	1	5506			
2	10025	1	5506			
2	10026	1	5506			
2	10027	1	5506			
2	10028	1	5506			
2	10029	1	5506			
2	10030	1	5506			
2	10031	1	5506			
2	10032	1	5520			
2	10033	1	5520			
2	10034	1	5520			
2	10035	1	5520			
2	10036	1	5520			
2	10037	1	5520			
2	10038	1	5520			
2	10039	1	5520			
2	10040	1	5520			
2	10041	1	5520			
2	10042	1	5520			
2	10043	1	5520			
2	10044	1	5520			
2	10045	1	5520			
2	10046	1	5520			
2	10047	1	5520			
2	10048	1	5520			
2	10049	1	5536			
2	10050	1	5536			
2	10051	1	5536			
2	10052	1	5536			
2	8511	1	332			
2	10053	1	5536			
2	10054	1	5536			
2	10055	1	5536			
2	10056	1	5536			
2	10057	1	5536			
2	8512	1	332			
2	10058	1	5536			
2	10059	1	5536			
2	10060	1	5536			
2	10063	1	5549			
2	10064	1	5549			
2	10065	1	5549			
2	10066	1	5549			
2	10067	1	5549			
2	10068	1	5549			
2	10069	1	5549			
2	10070	1	5555			
2	10071	1	5555			
2	10072	1	5555			
2	10073	1	5555			
2	10074	1	5555			
2	10075	1	5555			
2	10076	1	5555			
2	10077	1	5555			
2	10078	1	5562			
2	10079	1	5562			
2	10080	1	5562			
2	10081	1	5562			
2	10082	1	5562			
2	10083	1	5562			
2	10084	1	5562			
2	10085	1	5562			
2	10086	1	5562			
2	10087	1	5562			
2	10088	1	5562			
2	10089	1	5562			
2	10090	1	5573			
2	10091	1	5573			
2	10092	1	5573			
2	10093	1	5573			
2	10094	1	5573			
2	10095	1	5579			
2	10096	1	5579			
2	10097	1	5579			
2	10098	1	5579			
2	10099	1	5579			
2	10100	1	5579			
2	10101	1	5579			
2	10102	1	5595			
2	10103	1	5595			
2	10104	1	5595			
2	10105	1	5595			
2	10106	1	5595			
2	10107	1	5595			
2	10108	1	5595			
2	10109	1	5595			
2	10110	1	5595			
2	10111	1	5595			
2	10112	1	5595			
2	10113	1	5606			
2	10114	1	5606			
2	10115	1	5606			
2	10116	1	5606			
2	10117	1	5606			
2	10118	1	5606			
2	10119	1	5606			
2	10120	1	5606			
2	10121	1	5606			
2	10122	1	5606			
2	10123	1	5624			
2	10124	1	5624			
2	10125	1	5624			
2	10126	1	5624			
2	10127	1	5624			
2	10128	1	5624			
2	10129	1	5624			
2	10130	1	5624			
2	10131	1	5624			
2	10132	1	5624			
2	10133	1	5624			
2	10134	1	5634			
2	10135	1	5634			
2	10136	1	5634			
2	10137	1	5634			
2	10138	1	5634			
2	10139	1	5634			
2	10140	1	5634			
2	8218	1	137			
2	10172	1	5671			
2	10143	1	5655			
2	10144	1	5655			
2	10145	1	5655			
2	10146	1	5655			
2	10147	1	5655			
2	10148	1	5655			
2	10149	1	5655			
2	10150	1	5655			
2	10151	1	5655			
2	10152	1	5655			
2	10153	1	5655			
2	8531	1	341			
2	10154	1	5655			
2	10155	1	5655			
2	8870	1	588			
2	10156	1	5655			
2	8532	1	341			
2	10160	1	5671			
2	10161	1	5671			
2	10162	1	5671			
2	10163	1	5671			
3	1972	5	0	1	1146	
2	8533	1	341			
2	10164	1	5671			
2	10165	1	5671			
2	10166	1	5671			
2	8534	1	341			
2	10167	1	5671			
2	10168	1	5671			
2	10169	1	5671			
2	10170	1	5671			
2	8535	1	341			
2	10174	1	5684			
2	10175	1	5684			
2	10176	1	5684			
2	10177	1	5684			
2	8536	1	341			
2	10178	1	5684			
2	10181	1	5692			
2	10182	1	5692			
2	10183	1	5692			
2	8537	1	341			
2	10184	1	5696			
2	10185	1	5696			
2	10187	1	5700			
2	10188	1	5700			
2	10189	1	5700			
2	10190	1	5700			
2	10191	1	5703			
2	10192	1	5703			
2	10186	1	5696			
2	10194	1	5707			
2	10195	1	5707			
2	10196	1	5707			
2	10197	1	5711			
2	10198	1	5711			
2	10199	1	5711			
2	10200	1	5711			
2	10201	1	5736			
2	10202	1	5736			
2	10203	1	5739			
2	10204	1	5739			
2	10205	1	5742			
2	10206	1	5742			
2	10207	1	5745			
2	10208	1	5745			
2	10209	1	5756			
2	10210	1	5756			
2	10211	1	6025			
2	10212	1	6025			
2	10213	1	6028			
2	10214	1	6028			
2	10215	1	6045			
2	10171	1	5671			
2	10217	1	6080			
2	10218	1	6080			
2	10219	1	6091			
2	10220	1	6091			
2	10221	1	6108			
2	10222	1	6108			
2	10223	1	6117			
2	10224	1	6117			
2	8545	1	351			
2	10225	1	6140			
2	10227	1	6149			
2	10228	1	6149			
2	10229	1	6164			
2	10230	1	6164			
2	10231	1	6168			
2	10226	1	6140			
2	10233	1	6175			
2	10234	1	6175			
2	8547	1	351			
2	10235	1	6197			
2	10237	1	6200			
2	10232	1	6168			
2	10239	1	6203			
2	10236	1	6197			
2	10241	1	6206			
2	10238	1	6200			
2	10243	1	6397			
2	10244	1	6397			
2	10240	1	6203			
3	2054	7	0	2	136	1148	
2	10247	1	6415			
2	10248	1	6415			
2	10242	1	6206			
2	8550	1	351			
2	10245	1	6411			
3	2060	5	0	1	1150	
3	2061	5	0	1	1151	
2	10252	1	6427			
2	10253	1	6427			
2	10256	1	6441			
2	10257	1	6441			
2	10250	1	6419			
2	10251	1	6419			
2	10254	1	6437			
2	10261	1	6478			
2	10262	1	6478			
2	10263	1	6482			
2	10264	1	6482			
2	10265	1	6486			
2	10266	1	6486			
2	10267	1	6490			
2	10268	1	6490			
2	10269	1	6494			
2	10270	1	6494			
2	10271	1	6500			
2	10272	1	6500			
2	10273	1	6504			
2	10274	1	6504			
2	10275	1	6508			
2	10276	1	6508			
2	10277	1	6512			
2	10278	1	6512			
2	10279	1	6516			
2	10280	1	6516			
2	10281	1	6526			
2	10282	1	6526			
2	10283	1	6536			
2	10284	1	6536			
2	10285	1	6539			
2	10286	1	6539			
2	10287	1	6553			
2	10288	1	6553			
2	10289	1	6556			
2	8558	1	361			
2	10291	1	6566			
2	10292	1	6566			
2	10293	1	6569			
2	10294	1	6569			
2	8559	1	361			
2	10295	1	6572			
2	10296	1	6572			
2	10297	1	6575			
2	10298	1	6575			
2	10299	1	6580			
2	10300	1	6580			
2	10301	1	6584			
2	10302	1	6584			
2	10303	1	6587			
2	10304	1	6587			
2	10305	1	6592			
2	10307	1	6599			
2	10306	1	6592			
2	10309	1	6606			
2	10310	1	6606			
2	10311	1	6609			
2	10308	1	6599			
2	10313	1	6619			
2	10314	1	6619			
2	10315	1	6622			
2	10312	1	6609			
2	10317	1	6634			
2	10318	1	6634			
2	10319	1	6637			
2	8564	1	369			
2	10321	1	6792			
2	10320	1	6637			
2	10323	1	6795			
2	10193	1	5703			
2	10325	1	6817			
2	10326	1	6817			
2	10327	1	6817			
2	10328	1	6817			
2	10329	1	6817			
2	10330	1	6831			
2	10322	1	6792			
2	10332	1	6844			
2	10333	1	6844			
2	10334	1	6844			
2	10335	1	6844			
2	10336	1	6844			
2	10337	1	6857			
2	10331	1	6831			
2	10339	1	6866			
2	10340	1	6866			
2	10341	1	6866			
2	10342	1	6866			
2	10343	1	6866			
2	10344	1	6881			
2	10345	1	6881			
2	10346	1	6885			
2	10347	1	6885			
2	10348	1	6891			
2	10349	1	6891			
2	10350	1	6897			
2	10351	1	6897			
2	10352	1	6901			
2	10353	1	6901			
2	10354	1	6905			
2	10355	1	6905			
2	10356	1	6909			
2	9855	1	5264			
2	10357	1	6909			
2	10358	1	6916			
2	10360	1	6932			
2	10361	1	6932			
2	10362	1	6967			
2	10363	1	6967			
2	10364	1	6979			
2	10359	1	6916			
2	10365	1	6979			
2	10367	1	7003			
2	10368	1	7003			
2	10369	1	7006			
2	10370	1	7006			
2	10371	1	7023			
2	10372	1	7023			
2	10373	1	7023			
2	10374	1	7023			
2	8575	1	374			
2	10375	1	7028			
2	10377	1	7031			
2	10378	1	7031			
2	10379	1	7034			
2	10380	1	7034			
2	8576	1	374			
2	10381	1	7037			
2	10383	1	7041			
2	10382	1	7037			
2	10385	1	7049			
2	8577	1	374			
2	10386	1	7049			
2	10387	1	7049			
2	10389	1	7054			
2	10388	1	7049			
2	10391	1	7057			
2	10392	1	7057			
2	10393	1	7060			
2	10394	1	7060			
2	10395	1	7065			
2	10390	1	7054			
2	10397	1	7076			
2	10398	1	7076			
2	10399	1	7080			
2	10400	1	7080			
2	10401	1	7090			
2	10402	1	7090			
2	10403	1	7094			
2	10404	1	7094			
2	10405	1	7097			
2	10406	1	7097			
2	10407	1	7101			
2	10408	1	7101			
2	10409	1	7190			
2	10410	1	7190			
2	10411	1	7190			
2	10412	1	7190			
2	10413	1	7190			
2	10414	1	7198			
2	10415	1	7198			
2	10416	1	7198			
2	10417	1	7198			
2	10418	1	7198			
2	10419	1	7209			
2	10420	1	7209			
2	10421	1	7212			
2	10422	1	7212			
2	10423	1	7219			
2	10424	1	7219			
2	10425	1	7222			
2	10426	1	7222			
2	10427	1	7225			
2	10428	1	7225			
2	10429	1	7236			
2	10430	1	7236			
2	10431	1	7239			
2	10432	1	7239			
2	10433	1	7242			
2	10434	1	7242			
2	10435	1	7245			
2	10436	1	7245			
2	10437	1	7250			
2	10438	1	7250			
2	10439	1	7250			
2	10216	1	6045			
2	10440	1	7250			
2	10441	1	7250			
2	10443	1	7257			
2	10444	1	7257			
2	10445	1	7260			
2	10446	1	7260			
2	10447	1	7263			
2	10448	1	7263			
2	10449	1	7270			
2	10450	1	7270			
2	8590	1	389			
2	10451	1	7270			
2	10452	1	7270			
2	10454	1	7276			
2	10455	1	7276			
2	8591	1	389			
2	10456	1	7276			
2	10457	1	7276			
2	10459	1	7282			
2	10460	1	7282			
2	10461	1	7282			
2	10462	1	7282			
2	10463	1	7282			
2	10464	1	7288			
2	10465	1	7288			
2	10466	1	7288			
2	10467	1	7288			
2	10468	1	7288			
2	10469	1	7294			
2	10470	1	7294			
2	10471	1	7294			
2	10472	1	7294			
2	10473	1	7294			
2	10474	1	7301			
2	10475	1	7301			
2	10476	1	7304			
2	10477	1	7304			
2	10478	1	7304			
2	10479	1	7304			
2	10480	1	7304			
2	10481	1	7310			
2	10482	1	7310			
2	10483	1	7310			
2	10484	1	7310			
2	10485	1	7310			
2	10486	1	7402			
2	10487	1	7402			
2	10488	1	7409			
2	10489	1	7409			
2	10490	1	7412			
2	10491	1	7412			
2	10492	1	7421			
2	10493	1	7421			
2	10494	1	7489			
2	10495	1	7489			
2	10496	1	7531			
2	10497	1	7531			
2	10498	1	7531			
2	10499	1	7531			
2	10500	1	7531			
2	10501	1	7537			
2	10502	1	7537			
2	10503	1	7537			
2	10504	1	7537			
2	10505	1	7537			
2	10506	1	7543			
2	10507	1	7543			
2	10508	1	7543			
2	10509	1	7543			
2	10510	1	7543			
2	8602	1	400			
2	10511	1	7549			
2	10512	1	7549			
2	10513	1	7549			
2	10514	1	7549			
2	8603	1	400			
2	10516	1	7555			
2	10517	1	7555			
2	10518	1	7555			
2	10519	1	7555			
2	10521	1	7561			
2	10522	1	7561			
2	10523	1	7561			
2	10524	1	7561			
2	10525	1	7561			
2	10526	1	7567			
2	10527	1	7567			
2	10528	1	7567			
2	10529	1	7567			
2	10530	1	7567			
2	10531	1	7573			
2	10532	1	7573			
2	10533	1	7573			
2	10534	1	7573			
2	10535	1	7573			
2	10536	1	7579			
2	10537	1	7579			
2	10538	1	7582			
2	10539	1	7582			
2	10540	1	7589			
0	2349	7	1	2	9059	8716	
0	2350	3	1	2	9025	8717	
2	10541	1	7589			
2	10542	1	7592			
2	10543	1	7592			
2	10544	1	7595			
2	10545	1	7595			
2	10546	1	7712			
2	10547	1	7712			
2	10548	1	7715			
2	10549	1	7715			
2	10550	1	7724			
2	10551	1	7724			
2	10552	1	7762			
2	10553	1	7762			
2	10554	1	7765			
2	10555	1	7765			
2	10556	1	7772			
2	10557	1	7772			
2	10558	1	7775			
2	10559	1	7775			
2	10560	1	7778			
2	10561	1	7778			
2	10562	1	7800			
2	10563	1	7800			
2	10564	1	7803			
2	10565	1	7803			
2	10566	1	7812			
2	10567	1	7812			
2	10568	1	7826			
2	10569	1	7826			
2	8614	1	411			
2	10570	1	7829			
2	10571	1	7829			
2	10572	1	7836			
2	10573	1	7836			
2	8615	1	411			
2	10574	1	7839			
2	10515	1	7549			
2	10575	1	7839			
2	10576	1	7842			
2	10577	1	7842			
2	10578	1	7864			
2	10579	1	7864			
2	10580	1	7867			
2	10581	1	7867			
2	10582	1	7876			
2	10583	1	7876			
2	10584	1	7890			
2	10585	1	7890			
2	10246	1	6411			
2	10586	1	7893			
2	10587	1	7893			
2	10588	1	7900			
2	10589	1	7900			
2	10590	1	7903			
2	10591	1	7903			
2	10592	1	7906			
2	10593	1	7906			
2	10594	1	7932			
2	10595	1	7932			
2	10596	1	7935			
2	10597	1	7935			
2	10598	1	7940			
2	10599	1	7940			
2	10602	1	7957			
2	10600	1	7954			
2	10249	1	6415			
2	10603	1	7957			
2	10601	1	7954			
2	10608	1	7970			
2	10609	1	7970			
2	10606	1	7963			
2	10607	1	7963			
2	10610	1	7998			
2	10611	1	7998			
2	10612	1	8001			
2	10613	1	8001			
2	10614	1	8004			
2	10615	1	8004			
2	10616	1	8013			
2	10618	1	8017			
2	10620	1	8045			
2	10621	1	8045			
2	10622	1	8048			
2	10623	1	8048			
2	10619	1	8017			
2	10626	1	8064			
2	10624	1	8061			
2	10625	1	8061			
2	10627	1	8064			
2	10628	1	8079			
2	10630	1	8082			
2	10629	1	8079			
2	10631	1	8082			
2	10255	1	6437			
2	10636	1	8099			
2	10638	1	8102			
2	10639	1	8102			
2	10637	1	8099			
2	10179	1	5684			
2	8628	1	422			
2	10634	1	8096			
2	10635	1	8096			
2	8629	1	422			
2	10258	1	6441			
2	10259	1	6445			
2	10260	1	6445			
2	8640	1	435			
2	8641	1	435			
2	9870	1	5284			
2	9786	1	4425			
2	10180	1	5684			
2	8653	1	446			
3	2584	5	0	1	8754	
0	2585	7	1	3	8243	8769	8791	
0	2586	7	1	3	8245	8770	8792	
0	2587	7	1	3	8241	8771	8793	
0	2588	7	1	3	8239	8772	8794	
0	2589	7	1	3	8237	8773	8795	
3	2590	6	0	2	9077	140	
0	2591	7	1	3	8253	8774	8796	
0	2592	7	1	3	8235	8775	8797	
0	2593	7	1	3	8231	8776	8798	
0	2594	7	1	3	8227	8777	8799	
0	2595	7	1	3	8244	8813	8835	
0	2596	7	1	3	8246	8814	8836	
0	2597	7	1	3	8242	8815	8837	
0	2598	7	1	3	8240	8816	8838	
0	2599	7	1	3	8238	8817	8839	
0	2600	7	1	3	8254	8818	8840	
0	2601	7	1	3	8236	8819	8841	
0	2602	7	1	3	8232	8820	8842	
0	2603	7	1	3	8228	8821	8843	
0	2604	7	1	3	8194	8921	8943	
0	2605	7	1	3	8168	8899	8877	
0	2606	7	1	3	8195	8900	8878	
0	2607	7	1	3	8159	8901	8879	
0	2608	7	1	3	8192	8902	8880	
0	2609	7	1	3	8153	8903	8881	
0	2610	7	1	3	8151	8904	8882	
0	2611	7	1	3	8142	8905	8883	
0	2612	7	1	3	8140	8906	8884	
0	2613	7	1	3	8174	8907	8885	
0	2614	7	1	3	8170	8908	8886	
0	2615	7	1	3	8160	8922	8944	
0	2616	7	1	3	8193	8923	8945	
0	2617	7	1	3	8154	8924	8946	
0	2618	7	1	3	8152	8925	8947	
0	2619	7	1	3	8143	8926	8948	
0	2620	7	1	3	8141	8927	8949	
0	2621	7	1	3	8175	8928	8950	
0	2622	7	1	3	8171	8929	8951	
3	2623	5	0	1	9078	
0	2624	7	1	3	8198	9095	8872	
0	2625	7	1	2	8965	8994	
0	2626	7	1	3	8169	8930	8952	
0	2627	7	1	2	8966	8995	
0	2628	5	1	1	8642	
0	2629	5	1	1	8654	
0	2630	5	1	1	8666	
0	2631	5	1	1	8616	
0	2632	5	1	1	8630	
0	2633	5	1	1	8580	
0	2634	5	1	1	8592	
0	2635	5	1	1	8604	
0	2636	5	1	1	8565	
0	2637	5	1	1	8129	
0	2638	5	1	1	8643	
0	2639	5	1	1	8655	
0	2640	5	1	1	8667	
0	2641	5	1	1	8631	
0	2642	5	1	1	8581	
0	2643	5	1	1	8593	
0	2644	5	1	1	8605	
0	2645	5	1	1	8617	
0	2646	5	1	1	8566	
2	8210	1	137			
0	2653	5	10	1	8778	
0	2664	5	10	1	8800	
0	2681	5	10	1	8779	
0	2692	5	10	1	8801	
2	8676	1	468			
2	8677	1	468			
0	2703	7	1	3	8249	8780	8802	
0	2709	5	1	1	8678	
0	2710	5	1	1	8690	
0	2711	5	1	1	8704	
0	2712	5	1	1	8718	
0	2713	5	1	1	8726	
0	2714	5	1	1	8738	
0	2715	5	1	1	8161	
0	2716	5	1	1	8679	
0	2717	5	1	1	8705	
0	2718	5	1	1	8719	
0	2719	5	1	1	8727	
0	2720	5	1	1	8739	
0	2721	5	1	1	8691	
0	2728	5	10	1	8822	
0	2739	5	10	1	8844	
2	10316	1	6622			
2	8688	1	479			
0	2756	5	10	1	8823	
2	8689	1	479			
0	2767	5	10	1	8845	
0	2778	7	1	3	8250	8824	8846	
0	2779	5	10	1	8909	
0	2790	5	10	1	8887	
2	10324	1	6795			
2	8252	1	182			
0	2801	5	10	1	8931	
0	2812	5	10	1	8953	
0	2823	5	1	1	8278	
0	2824	5	1	1	8279	
0	2825	5	1	1	8289	
0	2826	5	1	1	8290	
0	2827	5	1	1	8300	
0	2828	5	1	1	8301	
0	2829	5	1	1	8311	
0	2830	5	1	1	8312	
0	2831	7	1	3	9060	8656	8280	
0	2832	7	1	3	9061	8668	8291	
0	2833	7	1	3	9062	8618	8302	
0	2834	7	1	3	9063	8632	8313	
0	2835	7	1	2	9026	8281	
0	2836	7	1	2	9027	8292	
0	2837	7	1	2	9028	8303	
0	2838	7	1	2	9029	8314	
0	2839	5	1	1	8406	
0	2840	5	1	1	8407	
0	2841	5	1	1	8417	
0	2842	5	1	1	8418	
0	2843	5	1	1	8428	
0	2844	5	1	1	8429	
0	2845	5	1	1	8439	
0	2846	5	1	1	8440	
0	2847	7	1	3	9064	8582	8408	
0	2848	7	1	3	9065	8594	8419	
0	2849	7	1	3	9066	8606	8430	
0	2850	7	1	3	9067	8567	8441	
0	2851	7	1	2	9030	8409	
0	2852	7	1	2	9031	8420	
0	2853	7	1	2	9032	8431	
0	2854	7	1	2	9033	8442	
0	2855	5	5	1	8513	
0	2861	5	5	1	8514	
2	10338	1	6857			
0	2867	7	1	2	292	8515	
0	2868	7	1	2	288	8516	
0	2869	7	1	2	280	8517	
0	2870	7	1	2	272	8518	
0	2871	7	1	2	264	8519	
0	2872	7	1	2	241	8520	
0	2873	7	1	2	233	8521	
0	2874	7	1	2	225	8522	
0	2875	7	1	2	217	8523	
0	2876	7	1	2	209	8524	
0	2882	5	8	1	8862	
2	8714	1	503			
2	8715	1	503			
0	2891	5	9	1	9079	
0	2901	5	1	1	8453	
0	2902	5	1	1	8462	
0	2903	5	1	1	8469	
0	2904	5	1	1	8470	
0	2905	5	1	1	8480	
0	2906	5	1	1	8481	
0	2907	7	1	2	8344	8463	
0	2908	7	1	3	8345	8680	8471	
0	2909	7	1	3	8346	8692	8482	
0	2910	7	1	2	8322	8454	
0	2911	7	1	2	8323	8472	
0	2912	7	1	2	8324	8483	
0	2913	5	1	1	8492	
0	2914	5	1	1	8493	
0	2915	5	1	1	8527	
0	2916	5	1	1	8528	
0	2917	5	1	1	8540	
0	2918	5	1	1	8541	
0	2919	7	1	3	9068	8706	8494	
0	2920	5	1	1	2349	
0	2921	7	1	3	9069	8728	8529	
0	2922	7	1	3	9070	8740	8542	
0	2923	7	1	2	9034	8495	
0	2924	7	1	2	9035	8530	
0	2925	7	1	2	9036	8543	
0	2926	5	1	1	8410	
0	2927	5	1	1	8411	
0	2928	5	1	1	8421	
0	2929	5	1	1	8422	
0	2930	5	1	1	8432	
0	2931	5	1	1	8433	
0	2932	5	1	1	8443	
0	2933	5	1	1	8444	
0	2934	7	1	3	8347	8583	8412	
0	2935	7	1	3	8348	8595	8423	
0	2936	7	1	3	8349	8607	8434	
0	2937	7	1	3	8350	8568	8445	
0	2938	7	1	2	8325	8413	
0	2939	7	1	2	8326	8424	
0	2940	7	1	2	8327	8435	
0	2941	7	1	2	8328	8446	
0	2942	5	5	1	8501	
2	8725	1	514			
0	2948	5	5	1	8502	
0	2954	7	1	2	372	8503	
0	2955	7	1	2	8561	8504	
0	2956	7	1	2	8552	8505	
0	2957	7	1	2	8539	8506	
0	2958	7	1	2	8526	8507	
0	2959	7	1	2	331	8508	
0	2960	7	1	2	323	8509	
0	2961	7	1	2	315	8510	
0	2962	7	1	2	307	8511	
0	2963	7	1	2	8460	8512	
0	2964	5	4	1	9084	
0	2969	7	1	2	8180	9085	
0	2970	7	1	2	86	9086	
0	2971	7	1	2	8182	9087	
0	2972	7	1	2	8183	9088	
0	2973	5	1	1	8496	
0	2974	5	1	1	8497	
0	2975	5	1	1	8531	
0	2976	5	1	1	8532	
0	2977	5	1	1	8544	
0	2978	5	1	1	8545	
0	2979	7	1	3	8351	8707	8498	
0	2980	7	1	2	8352	8720	
0	2981	7	1	3	8353	8729	8533	
0	2982	7	1	3	8354	8741	8546	
0	2983	7	1	2	8329	8499	
0	2984	3	1	2	8330	8721	
0	2985	7	1	2	8331	8534	
0	2986	7	1	2	8332	8547	
0	2987	5	1	1	8455	
0	2988	5	1	1	8464	
0	2989	5	1	1	8473	
0	2990	5	1	1	8474	
0	2991	5	1	1	8484	
0	2992	5	1	1	8485	
0	2993	7	1	2	8355	8465	
0	2994	7	1	3	8356	8681	8475	
0	2995	7	1	3	8357	8693	8486	
0	2996	7	1	2	8333	8456	
0	2997	7	1	2	8334	8476	
0	2998	7	1	2	8335	8487	
0	2999	5	1	1	8553	
2	8736	1	523			
2	8737	1	523			
2	10366	1	6979			
2	8260	1	194			
0	3006	5	1	1	8554	
0	3013	7	1	2	8358	8555	
0	3014	7	1	2	8359	8556	
0	3015	5	1	1	8282	
0	3016	5	1	1	8283	
0	3017	5	1	1	8293	
0	3018	5	1	1	8294	
0	3019	5	1	1	8304	
0	3020	5	1	1	8305	
0	3021	5	1	1	8315	
0	3022	5	1	1	8316	
0	3023	7	1	3	8360	8657	8284	
0	3024	7	1	3	8361	8669	8295	
0	3025	7	1	3	8362	8619	8306	
0	3026	7	1	3	8363	8633	8317	
0	3027	7	1	2	8336	8285	
0	3028	7	1	2	8337	8296	
0	3029	7	1	2	8338	8307	
0	3030	7	1	2	8339	8318	
0	3031	5	1	1	8557	
0	3032	5	1	1	8562	
0	3033	5	1	1	8535	
0	3034	5	1	1	8548	
0	3041	5	10	1	8910	
2	8747	1	534			
2	9890	1	5377			
0	3052	5	10	1	8888	
2	10376	1	7028			
2	8748	1	534			
2	8749	1	534			
0	3063	5	4	1	8996	
0	3068	5	2	1	8967	
0	3071	7	1	2	8188	8997	
0	3072	7	1	2	8186	8998	
0	3073	7	1	2	8189	8999	
0	3074	7	1	2	8187	9000	
0	3075	5	10	1	8932	
2	8754	1	549			
0	3086	5	10	1	8954	
2	10384	1	7041			
0	3097	5	10	1	8968	
2	8757	1	552			
0	3108	5	10	1	9001	
0	3119	5	10	1	8969	
0	3130	5	10	1	9002	
0	3141	5	1	1	8447	
0	3142	5	1	1	8450	
0	3143	5	1	1	8425	
0	3144	5	1	1	8436	
0	3145	5	1	1	8319	
0	3146	5	1	1	8414	
0	3147	5	10	1	8970	
2	8766	1	566			
2	8767	1	566			
2	10396	1	7065			
2	8768	1	566			
0	3158	5	10	1	9003	
0	3169	5	10	1	8971	
0	3180	5	10	1	9004	
2	9787	1	4425			
0	3194	5	1	1	8477	
0	3195	5	1	1	8488	
0	3196	5	1	1	8457	
0	3197	5	1	1	8466	
0	3198	5	1	1	8297	
0	3199	5	1	1	8308	
0	3203	5	1	1	8286	
2	8781	1	571			
2	8782	1	571			
2	8269	1	206			
2	8783	1	571			
2	8784	1	571			
2	8785	1	571			
2	8786	1	571			
2	8787	1	571			
2	8270	1	206			
2	8788	1	571			
2	9774	1	4418			
2	8789	1	571			
2	8790	1	571			
2	8271	1	206			
2	8806	1	574			
2	8807	1	574			
2	8808	1	574			
2	8809	1	574			
2	8810	1	574			
2	8811	1	574			
2	8812	1	574			
2	10442	1	7250			
0	3401	7	1	3	8658	9048	2824	
0	3402	7	1	3	8670	9049	2826	
0	3403	7	1	3	8620	9050	2828	
0	3404	7	1	3	8634	9051	2830	
0	3405	7	1	2	9037	2823	
0	3406	7	1	2	9038	2825	
0	3407	7	1	2	9039	2827	
0	3408	7	1	2	9040	2829	
0	3409	7	1	3	8584	9052	2840	
0	3410	7	1	3	8596	9053	2842	
0	3411	7	1	3	8608	9054	2844	
0	3412	7	1	3	8569	9055	2846	
0	3413	7	1	2	9041	2839	
0	3414	7	1	2	9042	2841	
0	3415	7	1	2	9043	2843	
0	3416	7	1	2	9044	2845	
2	10453	1	7270			
0	3444	7	1	2	8366	2902	
0	3445	7	1	3	8682	8367	2904	
0	3446	7	1	3	8694	8368	2906	
0	3447	7	1	2	8387	2901	
0	3448	7	1	2	8388	2903	
0	3449	7	1	2	8389	2905	
0	3450	7	1	3	8708	9056	2914	
0	3451	7	1	3	8730	9057	2916	
0	3452	7	1	3	8742	9058	2918	
0	3453	7	1	2	9045	2913	
0	3454	7	1	2	9046	2915	
0	3455	7	1	2	9047	2917	
0	3456	7	2	2	2920	2350	
0	3459	7	1	3	8585	8369	2927	
0	3460	7	1	3	8597	8370	2929	
0	3461	7	1	3	8609	8371	2931	
0	3462	7	1	3	8570	8372	2933	
0	3463	7	1	2	8390	2926	
0	3464	7	1	2	8391	2928	
0	3465	7	1	2	8392	2930	
0	3466	7	1	2	8393	2932	
2	10458	1	7276			
0	3481	7	1	3	8709	8373	2974	
0	3482	5	1	1	2980	
0	3483	7	1	3	8731	8374	2976	
0	3484	7	1	3	8743	8375	2978	
0	3485	7	1	2	8394	2973	
0	3486	7	1	2	8395	2975	
0	3487	7	1	2	8396	2977	
0	3488	7	1	2	8376	2988	
0	3489	7	1	3	8683	8377	2990	
0	3490	7	1	3	8695	8378	2992	
0	3491	7	1	2	8397	2987	
0	3492	7	1	2	8398	2989	
0	3493	7	1	2	8399	2991	
2	8834	1	577			
0	3502	7	1	2	8379	2999	
0	3503	7	1	2	8380	3006	
0	3504	7	1	3	8659	8381	3016	
0	3505	7	1	3	8671	8382	3018	
0	3506	7	1	3	8621	8383	3020	
0	3507	7	1	3	8635	8384	3022	
0	3508	7	1	2	8400	3015	
0	3509	7	1	2	8401	3017	
0	3510	7	1	2	8402	3019	
0	3511	7	1	2	8403	3021	
0	3512	6	1	2	8563	3031	
0	3513	6	1	2	8558	3032	
0	3514	6	1	2	8549	3033	
0	3515	6	1	2	8536	3034	
2	8220	1	137			
2	9797	1	4445			
0	3558	6	1	2	8451	3141	
0	3559	6	1	2	8448	3142	
0	3560	6	1	2	8437	3143	
0	3561	6	1	2	8426	3144	
0	3562	6	1	2	8415	3145	
0	3563	6	1	2	8320	3146	
0	3605	6	1	2	8489	3194	
0	3606	6	1	2	8478	3195	
0	3607	6	1	2	8467	3196	
0	3608	6	1	2	8458	3197	
0	3609	6	1	2	8309	3198	
0	3610	6	1	2	8298	3199	
2	8858	1	583			
2	8859	1	583			
3	3613	5	0	1	8461	
0	3614	7	1	2	9227	9235	
0	3615	7	1	2	8863	9236	
0	3616	7	1	3	8263	9097	8803	
0	3617	7	1	3	8265	9098	8804	
0	3618	7	1	3	8261	9099	8805	
0	3619	7	1	3	8259	9100	8806	
0	3620	7	1	3	8257	9101	8807	
0	3621	7	1	3	8251	9117	8808	
0	3622	7	1	3	8255	9118	8809	
0	3623	7	1	3	8233	9119	8810	
0	3624	7	1	3	8229	9120	8811	
0	3625	7	1	2	9228	9237	
0	3626	7	1	2	8864	9238	
0	3627	7	1	3	8264	9137	8847	
0	3628	7	1	3	8266	9138	8848	
0	3629	7	1	3	8262	9139	8849	
0	3630	7	1	3	8260	9140	8850	
0	3631	7	1	3	8258	9141	8851	
0	3632	7	1	3	8252	9157	8852	
0	3633	7	1	3	8256	9158	8853	
0	3634	7	1	3	8234	9159	8854	
0	3635	7	1	3	8230	9160	8855	
0	3636	7	1	2	9229	9239	
0	3637	7	1	2	8865	9240	
0	3638	7	1	3	8196	9284	8955	
0	3639	7	1	2	9230	9241	
0	3640	7	1	2	8866	9242	
0	3641	7	1	3	8136	9177	8889	
0	3642	7	1	3	8197	9258	8890	
0	3643	7	1	3	8157	9259	8891	
0	3644	7	1	3	8190	9260	8892	
0	3645	7	1	3	8184	9261	8893	
0	3646	7	1	3	8155	9262	8894	
0	3647	7	1	3	8178	9178	8895	
0	3648	7	1	3	8176	9179	8896	
0	3649	7	1	3	8172	9180	8897	
0	3650	7	1	3	8138	9181	8898	
0	3651	7	1	3	8158	9285	8956	
0	3652	7	1	3	8191	9286	8957	
0	3653	7	1	3	8185	9287	8958	
2	8286	1	210			
0	3654	7	1	3	8156	9288	8959	
0	3655	7	1	3	8179	9197	8960	
0	3656	7	1	3	8177	9198	8961	
0	3657	7	1	3	8173	9199	8962	
0	3658	7	1	3	8139	9200	8963	
0	3659	7	1	3	120	9324	9005	
0	3660	7	1	3	8137	9201	8964	
0	3661	7	1	3	118	9304	9006	
0	3662	7	1	3	8247	9121	8812	
0	3663	7	1	3	8248	9161	8856	
0	3664	3	1	2	2831	3401	
0	3665	3	1	2	2832	3402	
0	3666	3	1	2	2833	3403	
0	3667	3	1	2	2834	3404	
0	3668	3	1	3	2835	3405	8660	
0	3669	3	1	3	2836	3406	8672	
0	3670	3	1	3	2837	3407	8622	
0	3671	3	1	3	2838	3408	8636	
0	3672	3	1	2	2847	3409	
0	3673	3	1	2	2848	3410	
0	3674	3	1	2	2849	3411	
0	3675	3	1	2	2850	3412	
0	3676	3	1	3	2851	3413	8586	
0	3677	3	1	3	2852	3414	8598	
0	3678	3	1	3	2853	3415	8610	
0	3679	3	1	3	2854	3416	8571	
0	3680	7	1	2	8452	9217	
0	3681	7	1	2	8449	9218	
0	3682	7	1	2	8438	9219	
0	3683	7	1	2	8427	9220	
0	3684	7	1	2	8416	9221	
0	3685	7	1	2	8321	9222	
0	3686	7	1	2	8310	9223	
0	3687	7	1	2	8299	9224	
0	3688	7	1	2	8287	9225	
0	3689	7	1	2	8267	9226	
0	3691	5	8	1	9243	
2	8873	1	599			
2	8875	1	603			
2	8876	1	603			
0	3700	3	1	2	2907	3444	
0	3701	3	1	2	2908	3445	
0	3702	3	1	2	2909	3446	
0	3703	3	1	3	2911	3448	8684	
0	3704	3	1	3	2912	3449	8696	
0	3705	3	3	2	2910	3447	
0	3708	3	1	2	2919	3450	
0	3709	3	1	2	2921	3451	
0	3710	3	1	2	2922	3452	
0	3711	3	1	3	2923	3453	8710	
0	3712	3	1	3	2924	3454	8732	
0	3713	3	1	3	2925	3455	8744	
0	3715	3	1	2	2934	3459	
0	3716	3	1	2	2935	3460	
0	3717	3	1	2	2936	3461	
0	3718	3	1	2	2937	3462	
0	3719	3	1	3	2938	3463	8587	
0	3720	3	1	3	2939	3464	8599	
0	3721	3	1	3	2940	3465	8611	
0	3722	3	1	3	2941	3466	8572	
0	3723	7	1	2	8564	9244	
0	3724	7	1	2	8559	9245	
0	3725	7	1	2	8550	9246	
0	3726	7	1	2	8537	9247	
0	3727	7	1	2	8500	9249	
0	3728	7	1	2	8490	9250	
0	3729	7	1	2	8479	9251	
0	3730	7	1	2	8468	9252	
0	3731	7	1	2	8459	9253	
0	3732	3	8	2	9248	2958	
0	3738	7	1	2	8181	9254	
0	3739	7	1	2	87	9255	
0	3740	7	1	2	8149	9256	
0	3741	7	1	2	8150	9257	
0	3742	3	1	2	2979	3481	
0	3743	3	1	2	2981	3483	
0	3744	3	1	2	2982	3484	
0	3745	3	1	3	2983	3485	8711	
0	3746	3	1	3	2985	3486	8733	
0	3747	3	1	3	2986	3487	8745	
0	3748	3	1	2	2993	3488	
0	3749	3	1	2	2994	3489	
0	3750	3	1	2	2995	3490	
0	3751	3	1	3	2997	3492	8685	
0	3752	3	1	3	2998	3493	8697	
0	3753	5	1	1	8268	
0	3754	5	1	1	8269	
0	3755	5	1	1	8270	
0	3756	5	1	1	8271	
0	3757	3	1	2	3013	3502	
0	3758	7	1	3	8364	8644	8272	
0	3759	3	1	2	3014	3503	
0	3760	7	1	3	8365	8645	8273	
0	3761	7	1	2	8340	8274	
0	3762	7	1	2	8341	8275	
0	3763	3	1	2	3023	3504	
0	3764	3	1	2	3024	3505	
0	3765	3	1	2	3025	3506	
0	3766	3	1	2	3026	3507	
0	3767	3	1	3	3027	3508	8661	
0	3768	3	1	3	3028	3509	8673	
0	3769	3	1	3	3029	3510	8623	
0	3770	3	1	3	3030	3511	8637	
0	3771	6	3	2	3512	3513	
0	3775	6	3	2	3514	3515	
2	10520	1	7555			
0	3779	5	1	1	9089	
0	3780	5	1	1	9090	
0	3781	7	1	3	117	9305	9007	
0	3782	7	1	3	126	9306	9008	
0	3783	7	1	3	127	9307	9009	
0	3784	7	1	3	128	9308	9010	
0	3785	7	1	3	131	9325	9011	
0	3786	7	1	3	129	9326	9012	
0	3787	7	1	3	119	9327	9013	
0	3788	7	1	3	130	9328	9014	
0	3789	6	3	2	3558	3559	
0	3793	6	3	2	3560	3561	
0	3797	6	4	2	3562	3563	
0	3800	7	1	3	122	9344	9015	
0	3801	7	1	3	113	9345	9016	
0	3802	7	1	3	53	9346	9017	
0	3803	7	1	3	114	9347	9018	
0	3804	7	1	3	115	9348	9019	
0	3805	7	1	3	52	9364	9020	
0	3806	7	1	3	112	9365	9021	
0	3807	7	1	3	116	9366	9022	
0	3808	7	1	3	121	9367	9023	
0	3809	7	1	3	8199	9368	9024	
0	3810	6	2	2	3607	3608	
0	3813	6	2	2	3605	3606	
0	3816	7	2	2	3482	2984	
0	3819	3	2	2	2996	3491	
0	3822	5	1	1	8276	
0	3823	6	1	2	8277	3203	
0	3824	6	2	2	3609	3610	
0	3827	5	1	1	9384	
0	3828	3	1	2	3739	2970	
0	3829	3	1	2	3740	2971	
0	3830	3	1	2	3741	2972	
0	3831	3	1	2	3738	2969	
0	3834	5	1	1	3664	
0	3835	5	1	1	3665	
0	3836	5	1	1	3666	
0	3837	5	1	1	3667	
0	3838	5	1	1	3672	
0	3839	5	1	1	3673	
0	3840	5	1	1	3674	
0	3841	5	1	1	3675	
0	3842	3	9	2	3681	2868	
0	3849	3	8	2	3682	2869	
0	3855	3	8	2	3683	2870	
0	3861	3	8	2	3684	2871	
0	3867	3	8	2	3685	2872	
0	3873	3	10	2	3686	2873	
0	3881	3	8	2	3687	2874	
2	9775	1	4418			
0	3887	3	8	2	3688	2875	
0	3893	3	8	2	3689	2876	
0	3908	5	1	1	3701	
0	3909	5	1	1	3702	
0	3911	5	2	1	3700	
0	3914	5	1	1	3708	
0	3915	5	1	1	3709	
0	3916	5	1	1	3710	
0	3917	5	1	1	3715	
0	3918	5	1	1	3716	
0	3919	5	1	1	3717	
0	3920	5	1	1	3718	
0	3921	3	17	2	3724	2955	
2	8919	1	610			
2	8920	1	610			
0	3927	3	8	2	3725	2956	
0	3933	3	8	2	3726	2957	
0	3942	3	8	2	3727	2959	
2	8860	1	583			
0	3948	3	10	2	3728	2960	
0	3956	3	8	2	3729	2961	
0	3962	3	10	2	3730	2962	
0	3968	3	8	2	3731	2963	
0	3975	5	1	1	3742	
0	3976	5	1	1	3743	
0	3977	5	1	1	3744	
0	3978	5	1	1	3749	
0	3979	5	1	1	3750	
0	3980	7	1	3	8646	8385	3754	
0	3981	7	1	3	8647	8386	3756	
0	3982	7	1	2	8404	3753	
0	3983	7	1	2	8405	3755	
0	3984	5	2	1	3757	
0	3987	5	1	1	3759	
0	3988	5	1	1	3763	
0	3989	5	1	1	3764	
0	3990	5	1	1	3765	
0	3991	5	1	1	3766	
0	3998	7	1	3	9385	9329	9334	
0	4008	3	2	2	3723	2954	
0	4011	3	2	2	3680	2867	
0	4021	5	2	1	3748	
0	4024	6	1	2	8288	3822	
2	8941	1	613			
0	4027	5	1	1	9394	
2	8942	1	613			
0	4031	7	1	2	3828	9080	
0	4032	7	1	3	24	9231	9386	
0	4033	7	1	3	25	8867	9387	
0	4034	7	1	3	26	9232	9388	
0	4035	7	1	3	81	8868	9389	
0	4036	7	1	2	3829	9081	
0	4037	7	1	3	79	9233	9390	
0	4038	7	1	3	23	8869	9391	
0	4039	7	1	3	82	9234	9392	
0	4040	7	1	3	80	8870	9393	
0	4041	7	1	2	3830	9082	
0	4042	7	1	2	3831	9083	
0	4067	7	2	2	9397	8722	
0	4080	7	3	2	8723	9398	
0	4088	7	2	2	3834	3668	
0	4091	7	2	2	3835	3669	
0	4094	7	2	2	3836	3670	
0	4097	7	2	2	3837	3671	
0	4100	7	2	2	3838	3676	
0	4103	7	2	2	3839	3677	
0	4106	7	2	2	3840	3678	
0	4109	7	2	2	3841	3679	
0	4144	7	2	2	3908	3703	
0	4147	7	2	2	3909	3704	
0	4153	7	2	2	3914	3711	
0	4156	7	2	2	3915	3712	
0	4159	7	2	2	3916	3713	
2	9802	1	4456			
0	4183	3	1	2	3758	3980	
0	4184	3	1	2	3760	3981	
0	4185	3	1	3	3761	3982	8648	
0	4186	3	1	3	3762	3983	8649	
0	4188	5	2	1	9405	
0	4191	5	2	1	9408	
0	4196	7	1	3	9409	9406	9091	
0	4197	7	1	3	3987	9330	9335	
0	4198	7	1	2	3920	3722	
0	4199	5	1	1	9425	
0	4200	5	2	1	9411	
2	10604	1	7960			
0	4203	5	2	1	9414	
2	10605	1	7960			
2	8308	1	226			
0	4223	5	1	1	9421	
0	4224	5	1	1	9423	
0	4225	7	2	2	3918	3720	
0	4228	7	2	2	3919	3721	
2	9937	1	5424			
0	4231	7	2	2	3991	3770	
2	8309	1	226			
0	4234	7	2	2	3917	3719	
0	4237	7	2	2	3989	3768	
0	4240	7	2	2	3990	3769	
0	4243	7	2	2	3988	3767	
0	4246	7	2	2	3976	3746	
0	4249	7	2	2	3977	3747	
0	4252	7	2	2	3975	3745	
0	4255	7	2	2	3978	3751	
2	9938	1	5424			
0	4258	7	2	2	3979	3752	
2	8310	1	226			
0	4263	5	1	1	9427	
0	4264	6	2	2	4024	3823	
2	10617	1	8013			
0	4267	5	1	1	9429	
0	4268	7	1	2	8650	9498	
0	4269	5	1	1	9506	
0	4270	5	1	1	9585	
0	4271	7	1	2	9499	8651	
3	4272	5	0	1	4031	
0	4273	3	1	4	4032	4033	3614	3615	
0	4274	3	1	4	4034	4035	3625	3626	
3	4275	5	0	1	4036	
0	4276	3	1	4	4037	4038	3636	3637	
0	4277	3	1	4	4039	4040	3639	3640	
3	4278	5	0	1	4041	
3	4279	5	0	1	4042	
0	4280	7	3	2	9490	8662	
2	8991	1	619			
2	8992	1	619			
0	4284	7	5	2	9482	8674	
2	8993	1	619			
0	4290	7	7	2	8624	9472	
0	4297	7	1	2	9464	8638	
0	4298	7	2	2	9456	8588	
0	4301	7	3	2	9448	8600	
0	4305	7	4	2	9440	8612	
0	4310	7	5	2	9431	8573	
0	4316	7	3	2	8663	9491	
0	4320	7	4	2	8675	9483	
0	4325	7	6	2	8625	9473	
0	4331	7	1	2	8639	9465	
0	4332	7	3	2	8589	9457	
0	4336	7	5	2	8601	9449	
2	10632	1	8093			
0	4342	7	6	2	8613	9441	
2	10633	1	8093			
0	4349	7	8	2	8574	9432	
0	4357	5	8	1	9577	
0	4364	5	12	1	9567	
0	4379	7	5	2	9559	8686	
0	4385	7	7	2	8698	9549	
0	4392	7	1	2	9541	8712	
0	4396	7	3	2	9533	8734	
0	4400	7	4	2	9525	8746	
0	4405	5	7	1	9508	
0	4418	5	8	1	9578	
0	4425	5	12	1	9568	
2	9023	1	625			
0	4440	7	4	2	8687	9560	
2	9024	1	625			
0	4445	7	6	2	8699	9550	
0	4451	7	1	2	8713	9542	
2	9946	1	5431			
0	4456	7	5	2	8735	9534	
0	4462	7	6	2	8747	9526	
0	4477	5	8	1	9509	
2	9947	1	5431			
2	9948	1	5431			
0	4515	5	1	1	4183	
0	4516	5	1	1	4184	
2	9039	1	1080			
0	4521	5	1	1	9587	
0	4523	5	1	1	9589	
0	4524	5	3	1	4198	
0	4532	5	3	1	9586	
0	4547	7	1	3	9507	9369	9374	
0	4575	4	2	2	8626	9474	
0	4605	4	2	2	8627	9475	
0	4608	4	2	2	8575	9433	
0	4627	4	2	2	8700	9551	
0	4646	4	2	2	8701	9552	
2	9073	1	1157			
2	9074	1	1219			
2	9075	1	1219			
0	4701	6	1	2	9424	4223	
0	4702	6	1	2	9422	4224	
2	9076	1	1219			
0	4720	5	1	1	9591	
0	4721	6	1	2	9592	4263	
0	4724	5	1	1	9616	
0	4725	5	1	1	9614	
0	4726	5	1	1	9622	
0	4727	5	1	1	9620	
0	4728	5	1	1	9618	
0	4729	5	1	1	9604	
0	4730	5	1	1	9602	
0	4731	5	1	1	9600	
0	4732	5	1	1	9598	
0	4733	5	1	1	9612	
2	9082	1	1583			
0	4734	5	1	1	9610	
0	4735	5	1	1	9608	
3	4737	7	0	2	4273	8223	
3	4738	7	0	2	4274	8224	
3	4739	7	0	2	4276	8225	
3	4740	7	0	2	4277	8226	
0	4736	5	1	1	9606	
0	4741	7	1	3	9395	9096	9093	
2	9092	1	1660			
2	9093	1	1755			
2	9156	1	2739			
0	4855	5	1	1	9399	
0	4856	6	1	2	9400	2712	
2	9106	1	2653			
2	9116	1	2664			
0	4908	6	1	2	9401	2718	
0	4909	5	1	1	9402	
2	10290	1	6556			
0	4939	7	3	2	4515	4185	
0	4942	7	1	2	4516	4186	
0	4947	5	1	1	9403	
0	4953	7	1	3	9624	9410	3779	
0	4954	7	1	3	9407	9626	3780	
0	4955	7	1	3	9627	9625	9092	
0	4956	7	1	3	9613	9309	9314	
0	4957	7	1	3	9611	9310	9315	
0	4958	7	1	3	9609	9311	9316	
0	4959	7	1	3	9607	9312	9317	
0	4960	7	1	3	9623	9331	9336	
0	4961	7	1	3	9621	9332	9337	
2	9126	1	2681			
0	4965	5	1	1	9632	
0	4966	5	1	1	9634	
0	4967	5	1	1	9636	
0	4968	5	1	1	9638	
0	4972	5	1	1	9646	
0	4973	5	1	1	9648	
0	4974	5	1	1	9650	
0	4975	6	1	2	9651	4199	
0	4976	5	1	1	9417	
0	4977	5	1	1	9418	
0	4978	7	1	3	9415	9412	9419	
0	4979	7	1	3	9630	9628	9420	
0	4980	7	1	3	9605	9349	9354	
0	4981	7	1	3	9603	9350	9355	
0	4982	7	1	3	9601	9351	9356	
0	4983	7	1	3	9599	9352	9357	
0	4984	7	1	3	9619	9370	9375	
0	4985	7	1	3	9617	9371	9376	
0	4986	7	1	3	9615	9372	9377	
0	4987	7	1	3	9396	9373	9378	
2	8990	1	619			
2	8665	1	457			
2	9136	1	2692			
0	5049	6	2	2	4701	4702	
2	9145	1	2728			
0	5052	5	1	1	9640	
0	5053	5	1	1	9642	
0	5054	5	1	1	9644	
0	5055	5	1	1	9652	
0	5056	5	1	1	9654	
0	5057	6	1	2	9428	4720	
0	5058	5	1	1	9656	
0	5059	6	1	2	9657	4267	
0	5060	7	1	4	4724	4725	4269	4027	
0	5061	7	1	4	4726	4727	3827	4728	
0	5062	7	1	4	4729	4730	4731	4732	
0	5063	7	1	4	4733	4734	4735	4736	
2	9146	1	2728			
0	5065	7	1	2	9722	9569	
0	5066	7	1	3	9730	9723	9742	
0	5067	7	1	2	9768	9570	
0	5068	7	1	3	9776	9769	9788	
0	5069	5	1	1	9500	
0	5070	6	1	2	9501	2628	
0	5071	5	1	1	9492	
0	5072	6	1	2	9493	2629	
0	5073	5	1	1	9484	
0	5074	6	1	2	9485	2630	
0	5075	5	1	1	9476	
0	5076	6	1	2	9477	2631	
0	5077	5	1	1	9466	
0	5078	6	1	2	9467	2632	
0	5079	5	1	1	9458	
0	5080	6	1	2	9459	2633	
0	5081	5	1	1	9450	
0	5082	6	1	2	9451	2634	
0	5083	5	1	1	9442	
0	5084	6	1	2	9443	2635	
0	5085	5	1	1	9434	
0	5086	6	1	2	9435	2636	
0	5087	5	1	1	9823	
0	5088	6	1	2	9502	2638	
0	5089	5	1	1	9503	
0	5090	6	1	2	9494	2639	
0	5091	5	1	1	9495	
0	5092	6	1	2	9486	2640	
0	5093	5	1	1	9487	
0	5094	6	1	2	9468	2641	
0	5095	5	1	1	9469	
0	5096	6	1	2	9460	2642	
0	5097	5	1	1	9461	
0	5098	6	1	2	9452	2643	
0	5099	5	1	1	9453	
0	5100	6	1	2	9444	2644	
0	5101	5	1	1	9445	
0	5102	6	1	2	9478	2645	
0	5103	5	1	1	9479	
0	5104	6	1	2	9436	2646	
0	5105	5	1	1	9437	
0	5106	5	1	1	9561	
0	5107	6	1	2	9562	2709	
0	5108	5	1	1	9553	
0	5109	6	1	2	9554	2710	
0	5110	5	1	1	9543	
0	5111	6	1	2	9544	2711	
0	5112	6	1	2	8724	4855	
0	5113	5	1	1	9535	
0	5114	6	1	2	9536	2713	
0	5115	5	1	1	9527	
0	5116	6	1	2	9528	2714	
0	5117	7	1	2	9731	9743	
0	5118	7	1	2	9732	9744	
0	5119	7	1	2	8162	9761	
0	5120	5	1	1	9829	
0	5121	6	1	2	9563	2716	
0	5122	5	1	1	9564	
0	5123	6	1	2	9545	2717	
0	5124	5	1	1	9546	
0	5125	6	1	2	8725	4909	
0	5126	6	1	2	9537	2719	
0	5127	5	1	1	9538	
0	5128	6	1	2	9529	2720	
0	5129	5	1	1	9530	
0	5130	6	1	2	9555	2721	
0	5131	5	1	1	9556	
0	5132	7	1	2	9777	9789	
0	5133	7	1	2	9778	9790	
0	5135	5	1	1	9531	
0	5136	5	1	1	9539	
0	5137	6	1	2	9510	4521	
0	5138	5	1	1	9511	
0	5139	5	1	1	9547	
0	5140	6	1	2	9548	4947	
0	5141	5	1	1	9480	
0	5142	5	1	1	9470	
0	5143	5	1	1	9496	
0	5144	5	1	1	9488	
0	5145	6	1	2	9504	4523	
0	5146	5	1	1	9505	
0	5147	4	1	2	4953	4196	
0	5148	4	1	2	4954	4955	
2	8214	1	137			
0	5150	5	2	1	9817	
0	5153	6	1	2	9635	4965	
0	5154	6	1	2	9633	4966	
0	5155	6	1	2	9639	4967	
0	5156	6	1	2	9637	4968	
0	5157	5	2	1	9820	
2	9166	1	2756			
0	5160	6	1	2	9649	4972	
0	5161	6	1	2	9647	4973	
0	5162	6	1	2	9426	4974	
0	5163	7	1	3	9629	9416	4976	
0	5164	7	1	3	9413	9631	4977	
0	5165	7	1	3	4942	9353	9358	
0	5166	5	2	1	9579	
0	5172	5	1	1	9825	
0	5176	5	1	1	9827	
2	8833	1	577			
0	5198	5	1	1	9831	
2	9175	1	2767			
2	9176	1	2767			
0	5223	5	1	1	9565	
0	5224	5	1	1	9557	
0	5225	5	1	1	9580	
0	5226	5	1	1	9571	
0	5227	5	1	1	9446	
0	5228	5	1	1	9438	
0	5229	5	1	1	9462	
0	5230	5	1	1	9454	
0	5232	6	1	2	9643	5052	
0	5233	6	1	2	9641	5053	
0	5234	6	1	2	9655	5055	
0	5235	6	1	2	9653	5056	
0	5236	6	2	2	4721	5057	
0	5239	6	1	2	9430	5058	
3	5240	7	0	3	5060	5061	4270	
0	5241	5	1	1	9833	
0	5242	6	1	2	8652	5069	
0	5243	6	1	2	8664	5071	
0	5244	6	1	2	8676	5073	
0	5245	6	1	2	8628	5075	
0	5246	6	1	2	8640	5077	
0	5247	6	1	2	8590	5079	
0	5248	6	1	2	8602	5081	
0	5249	6	1	2	8614	5083	
0	5250	6	1	2	8576	5085	
0	5252	6	1	2	8653	5089	
0	5253	6	1	2	8665	5091	
0	5254	6	1	2	8677	5093	
0	5255	6	1	2	8641	5095	
0	5256	6	1	2	8591	5097	
0	5257	6	1	2	8603	5099	
0	5258	6	1	2	8615	5101	
0	5259	6	1	2	8629	5103	
0	5260	6	1	2	8577	5105	
0	5261	6	1	2	8688	5106	
0	5262	6	1	2	8702	5108	
0	5263	6	1	2	8714	5110	
0	5264	6	10	2	5112	4856	
2	9186	1	2779			
0	5274	6	1	2	8736	5113	
0	5275	6	1	2	8748	5115	
0	5282	6	1	2	8689	5122	
0	5283	6	1	2	8715	5124	
0	5284	6	15	2	4908	5125	
0	5298	6	1	2	8737	5127	
0	5299	6	1	2	8749	5129	
0	5300	6	1	2	8703	5131	
2	9194	1	2790			
0	5303	6	1	2	9540	5135	
0	5304	6	1	2	9532	5136	
0	5305	6	1	2	9588	5138	
0	5306	6	1	2	9404	5139	
0	5307	6	1	2	9471	5141	
0	5308	6	1	2	9481	5142	
0	5309	6	1	2	9489	5143	
0	5310	6	1	2	9497	5144	
0	5311	6	1	2	9590	5146	
0	5312	5	1	1	9836	
2	9196	1	2790			
0	5315	6	3	2	5153	5154	
0	5319	6	4	2	5155	5156	
0	5324	6	3	2	5160	5161	
0	5328	6	4	2	5162	4975	
0	5331	4	1	2	5163	4978	
0	5332	4	1	2	5164	4979	
0	5346	3	2	2	9512	5119	
2	9206	1	2801			
0	5363	6	1	2	9558	5223	
0	5364	6	1	2	9566	5224	
0	5365	6	1	2	9572	5225	
0	5366	6	1	2	9581	5226	
0	5367	6	1	2	9439	5227	
0	5368	6	1	2	9447	5228	
0	5369	6	1	2	9455	5229	
0	5370	6	1	2	9463	5230	
0	5371	6	2	2	5148	5147	
0	5377	6	2	2	5232	5233	
0	5382	6	2	2	5234	5235	
0	5385	6	2	2	5239	5059	
3	5388	7	0	3	5062	5063	5241	
0	5389	6	8	2	5242	5070	
0	5396	6	12	2	5243	5072	
0	5407	6	12	2	5244	5074	
2	9216	1	2812			
0	5418	6	5	2	5245	5076	
0	5424	6	7	2	5246	5078	
0	5431	6	10	2	5247	5080	
0	5441	6	11	2	5248	5082	
0	5452	6	10	2	5249	5084	
0	5462	6	7	2	5250	5086	
0	5469	5	1	1	9666	
0	5470	6	8	2	5088	5252	
0	5477	6	12	2	5090	5253	
0	5488	6	11	2	5092	5254	
0	5498	6	9	2	5094	5255	
2	9234	1	2882			
0	5506	6	15	2	5096	5256	
0	5520	6	17	2	5098	5257	
0	5536	6	14	2	5100	5258	
0	5549	6	7	2	5102	5259	
0	5555	6	8	2	5104	5260	
0	5562	6	12	2	5261	5107	
0	5573	6	5	2	5262	5109	
0	5579	6	7	2	5263	5111	
0	5595	6	11	2	5274	5114	
0	5606	6	10	2	5275	5116	
0	5616	6	1	2	9762	2715	
0	5617	5	1	1	9763	
0	5618	5	1	1	9724	
0	5619	5	1	1	9725	
0	5620	5	1	1	9733	
0	5621	5	1	1	9734	
0	5622	5	1	1	9747	
0	5624	6	11	2	5121	5282	
0	5634	6	9	2	5123	5283	
0	5655	6	17	2	5126	5298	
2	9267	1	3041			
0	5671	6	14	2	5128	5299	
0	5684	6	7	2	5130	5300	
0	5690	5	1	1	9779	
0	5691	5	1	1	9780	
0	5692	6	3	2	5303	5304	
2	9995	1	5477			
2	8367	1	251			
0	5696	6	3	2	5137	5305	
0	5700	6	4	2	5306	5140	
0	5703	6	3	2	5307	5308	
0	5707	6	3	2	5309	5310	
0	5711	6	4	2	5145	5311	
2	9996	1	5477			
2	8368	1	251			
2	9279	1	3063			
0	5726	7	1	2	9842	9582	
0	5727	5	1	1	9694	
0	5728	5	1	1	9714	
0	5730	5	1	1	9770	
0	5731	5	1	1	9792	
0	5732	5	1	1	9771	
0	5733	5	1	1	9809	
0	5734	5	1	1	9513	
0	5735	5	1	1	9810	
0	5736	6	2	2	5365	5366	
2	9280	1	3063			
2	9281	1	3063			
0	5739	6	2	2	5363	5364	
0	5742	6	2	2	5369	5370	
0	5745	6	2	2	5367	5368	
0	5755	5	1	1	9844	
0	5756	6	2	2	5332	5331	
2	8215	1	137			
2	9292	1	3075			
2	9293	1	3075			
2	9302	1	3086			
2	10141	1	5634			
2	9303	1	3086			
2	9313	1	3097			
2	9321	1	3108			
2	9322	1	3108			
2	9323	1	3108			
2	8703	1	490			
0	5954	7	1	2	9846	9754	
0	5955	6	1	2	8163	5617	
0	5956	5	1	1	9885	
2	10006	1	5488			
2	10142	1	5634			
2	9329	1	3119			
2	9330	1	3119			
2	9331	1	3119			
2	9332	1	3119			
2	9333	1	3119			
2	9334	1	3130			
0	6005	7	1	2	9856	9798	
0	6006	7	1	2	9857	9799	
2	9335	1	3130			
2	9336	1	3130			
2	9337	1	3130			
2	9338	1	3130			
0	6023	5	1	1	9887	
0	6024	6	1	2	9888	5312	
0	6025	5	2	1	9871	
2	9339	1	3130			
0	6028	5	2	1	9878	
2	9340	1	3130			
2	9341	1	3130			
2	9342	1	3130			
0	6044	5	1	1	9893	
0	6045	3	2	2	9843	5726	
2	9343	1	3130			
0	6065	5	1	1	9834	
0	6066	6	1	2	9835	5054	
0	6067	5	1	1	9889	
0	6068	5	1	1	9891	
0	6069	6	1	2	9892	5755	
0	6071	7	1	2	9977	9687	
0	6072	7	1	3	9985	9978	9690	
0	6073	7	1	4	9997	9979	9695	9986	
0	6074	7	1	4	10078	9726	9748	9735	
0	6075	7	1	2	9895	9658	
0	6076	7	1	3	9903	9896	9661	
0	6077	7	1	4	9915	9897	9667	9904	
0	6078	7	1	4	10123	9772	9793	9781	
0	6079	5	1	1	9927	
0	6080	7	2	4	9905	9928	9916	9898	
2	9359	1	3158			
0	6083	7	1	2	9906	9662	
0	6084	7	1	3	9917	9668	9907	
0	6085	7	1	3	9929	9918	9908	
0	6086	7	1	2	9909	9663	
0	6087	7	1	3	9669	9919	9910	
0	6088	7	1	2	9920	9670	
0	6089	7	1	2	9930	9921	
0	6090	7	1	2	9922	9671	
0	6091	7	2	5	9939	9970	9949	9932	9960	
0	6094	7	1	2	9933	9673	
0	6095	7	1	3	9940	9934	9675	
0	6096	7	1	4	9950	9935	9678	9941	
0	6097	7	1	5	9961	9951	9936	9682	9942	
2	9353	1	3147			
0	6098	7	1	2	9943	9676	
0	6099	7	1	3	9952	9679	9944	
0	6100	7	1	4	9962	9953	9683	9945	
0	6101	7	1	5	8130	9971	9954	9963	9946	
0	6102	7	1	2	9680	9955	
0	6103	7	1	3	9964	9956	9684	
0	6104	7	1	4	8131	9972	9957	9965	
0	6105	7	1	2	9966	9685	
0	6106	7	1	3	8132	9973	9967	
0	6107	7	1	2	8133	9974	
0	6108	7	2	4	10063	9998	9987	9980	
0	6111	7	1	2	9988	9691	
0	6112	7	1	3	9999	9696	9989	
0	6113	7	1	3	10064	10000	9990	
0	6114	7	1	2	9991	9692	
0	6115	7	1	3	10001	9697	9992	
0	6116	7	1	2	10002	9698	
0	6117	7	2	5	10070	10049	10032	10017	10008	
0	6120	7	1	2	10009	9700	
0	6121	7	1	3	10018	10010	9703	
0	6122	7	1	4	10033	10011	9708	10019	
0	6123	7	1	5	10050	10034	10012	9715	10020	
0	6124	7	1	2	10021	9704	
0	6125	7	1	3	10035	9709	10022	
0	6126	7	1	4	10051	10036	9716	10023	
0	6127	7	1	4	10071	10037	10024	10052	
0	6128	7	1	2	10025	9705	
0	6129	7	1	3	10038	9710	10026	
0	6130	7	1	4	10053	10039	9717	10027	
0	6131	7	1	2	10040	9711	
0	6132	7	1	3	10054	10041	9718	
0	6133	7	1	3	10072	10042	10055	
0	6134	7	1	2	10043	9712	
0	6135	7	1	3	10056	10044	9719	
0	6136	7	1	2	10057	9720	
0	6137	7	1	2	10065	10003	
0	6138	7	1	2	10073	10058	
0	6139	5	1	1	10090	
0	6140	7	2	4	9736	10091	10079	9727	
2	9360	1	3158			
2	9361	1	3158			
0	6143	7	1	3	10080	9749	9737	
0	6144	7	1	3	10092	10081	9738	
0	6145	7	1	3	9750	10082	9739	
0	6146	7	1	2	10083	9751	
0	6147	7	1	2	10093	10084	
0	6148	7	1	2	10085	9752	
0	6149	7	2	5	9847	9764	10102	10095	10113	
2	9362	1	3158			
2	9363	1	3158			
0	6152	7	1	2	10096	9593	
0	6153	7	1	3	9848	10097	9755	
0	6154	7	1	4	10103	10098	9757	9849	
0	6155	7	1	5	10114	10104	10099	9514	9850	
0	6156	7	1	3	10105	9758	9851	
0	6157	7	1	4	10115	10106	9515	9852	
0	6158	7	1	5	8164	9765	10107	10116	9853	
0	6159	7	1	2	9759	10108	
0	6160	7	1	3	10117	10109	9516	
0	6161	7	1	4	8165	9766	10110	10118	
0	6162	7	1	2	10119	9517	
0	6163	7	1	3	8166	9767	10120	
0	6164	6	2	2	5616	5955	
0	6168	7	2	4	10174	10124	9782	9773	
0	6171	7	1	3	10125	9794	9783	
0	6172	7	1	3	10175	10126	9784	
0	6173	7	1	3	10127	9795	9785	
0	6174	7	1	2	10128	9796	
0	6175	7	2	5	9811	10160	10143	9858	10134	
0	6178	7	1	2	10135	9595	
0	6179	7	1	3	9859	10136	9800	
0	6180	7	1	4	10144	10137	9803	9860	
0	6181	7	1	5	10161	10145	10138	9518	9861	
0	6182	7	1	3	10146	9804	9862	
0	6183	7	1	4	10162	10147	9519	9863	
0	6184	7	1	4	9812	10148	9864	10163	
0	6185	7	1	3	10149	9805	9865	
0	6186	7	1	4	10164	10150	9520	9866	
0	6187	7	1	2	10151	9806	
0	6188	7	1	3	10165	10152	9521	
0	6189	7	1	3	9813	10153	10166	
0	6190	7	1	2	10154	9807	
0	6191	7	1	3	10167	10155	9522	
0	6192	7	1	2	10168	9523	
0	6193	7	1	2	10176	10129	
0	6194	7	1	2	9814	10169	
2	10015	1	5498			
0	6197	5	2	1	10181	
0	6200	5	2	1	10184	
0	6203	5	2	1	10191	
0	6206	5	2	1	10194	
2	10016	1	5498			
0	6221	6	1	2	9837	6023	
0	6234	5	1	1	10209	
0	6235	6	1	2	10210	6044	
2	9396	1	3705			
2	8256	1	188			
2	9404	1	3732			
0	6373	5	1	1	10201	
0	6374	5	1	1	10203	
0	6375	5	1	1	10205	
0	6376	5	1	1	10207	
0	6377	6	1	2	9645	6065	
0	6378	6	1	2	9845	6068	
0	6382	3	1	4	4268	6071	6072	6073	
0	6386	3	1	4	9583	5065	5066	6074	
0	6388	3	1	4	4271	6075	6076	6077	
0	6392	3	1	4	9584	5067	5068	6078	
2	9412	1	3789			
2	8216	1	137			
0	6397	3	2	5	4297	6094	6095	6096	6097	
2	9413	1	3789			
0	6411	3	2	2	9693	6116	
2	9416	1	3793			
0	6415	3	3	5	4331	6120	6121	6122	6123	
0	6419	3	2	2	9713	6136	
0	6427	3	2	5	4392	6152	6153	6154	6155	
0	6434	5	1	1	9854	
2	9420	1	3797			
0	6437	3	2	2	9791	6174	
0	6441	3	3	5	4451	6178	6179	6180	6181	
0	6445	3	2	2	9808	6192	
2	8219	1	137			
0	6448	5	1	1	9867	
0	6449	5	1	1	9868	
2	9426	1	3816			
3	6466	6	0	2	6221	6024	
0	6469	5	1	1	9874	
0	6470	5	1	1	9875	
0	6471	5	1	1	9881	
0	6472	5	1	1	9882	
0	6473	7	1	3	9872	9818	9876	
0	6474	7	1	3	10211	9838	9877	
0	6475	7	1	3	9879	9821	9883	
0	6476	7	1	3	10213	9840	9884	
0	6477	6	1	2	9894	6234	
0	6478	6	2	2	10215	8200	
0	6482	3	2	4	9659	6083	6084	6085	
0	6486	4	2	3	9660	6086	6087	
0	6490	3	2	3	9664	6088	6089	
0	6494	4	2	2	9665	6090	
0	6500	3	2	5	9674	6098	6099	6100	6101	
0	6504	3	2	4	9677	6102	6103	6104	
0	6508	3	2	3	9681	6105	6106	
0	6512	3	2	2	9686	6107	
0	6516	3	2	4	9688	6111	6112	6113	
0	6526	4	2	3	9689	6114	6115	
0	6536	3	2	4	9706	6131	6132	6133	
0	6539	3	2	5	9701	6124	6125	6126	6127	
0	6553	4	2	3	9707	6134	6135	
0	6556	4	2	4	9702	6128	6129	6130	
0	6566	3	2	4	9573	5117	6143	6144	
0	6569	4	2	3	9574	5118	6145	
0	6572	3	2	3	9745	6146	6147	
0	6575	4	2	2	9746	6148	
2	8258	1	191			
0	6580	3	2	5	9594	5954	6156	6157	6158	
0	6584	3	2	4	9756	6159	6160	6161	
0	6587	3	2	3	9760	6162	6163	
0	6592	3	2	4	9575	5132	6171	6172	
0	6599	4	2	3	9576	5133	6173	
0	6606	3	2	4	9801	6187	6188	6189	
0	6609	3	2	5	9596	6005	6182	6183	6184	
0	6619	4	2	3	9802	6190	6191	
0	6622	4	2	4	9597	6006	6185	6186	
0	6630	6	1	2	10204	6373	
0	6631	6	1	2	10202	6374	
0	6632	6	1	2	10208	6375	
0	6633	6	1	2	10206	6376	
0	6634	6	2	2	6377	6066	
0	6637	6	2	2	6069	6378	
0	6640	5	1	1	10229	
3	6641	7	0	2	10221	10223	
3	6643	7	0	2	10225	10227	
3	6646	7	0	2	10231	10233	
2	8221	1	137			
3	6648	7	0	2	10217	10219	
0	6650	6	1	2	9975	2637	
2	9463	1	3861			
0	6651	5	1	1	9976	
0	6653	5	1	1	9899	
0	6655	5	1	1	9900	
0	6657	5	1	1	9911	
0	6659	5	1	1	9912	
0	6660	6	1	2	9923	5087	
0	6661	5	1	1	9924	
0	6662	6	1	2	9925	5469	
0	6663	5	1	1	9926	
0	6664	7	1	2	10220	8134	
0	6666	5	1	1	9937	
0	6668	5	1	1	9947	
0	6670	5	1	1	9958	
0	6672	5	1	1	9968	
0	6675	5	1	1	10224	
0	6680	5	1	1	9993	
0	6681	5	1	1	9994	
0	6682	5	1	1	10028	
0	6683	5	1	1	10029	
0	6689	6	1	2	10086	5120	
0	6690	5	1	1	10087	
0	6691	6	1	2	10088	5622	
0	6692	5	1	1	10089	
0	6693	7	1	2	10228	8167	
0	6695	5	1	1	10100	
0	6698	5	1	1	10111	
0	6699	6	1	2	10121	5956	
0	6700	5	1	1	10122	
0	6703	5	1	1	10234	
0	6708	5	1	1	10187	
0	6709	5	1	1	10188	
0	6710	5	1	1	10197	
0	6711	5	1	1	10198	
0	6712	7	1	3	10185	10182	10189	
0	6713	7	1	3	10237	10235	10190	
0	6714	7	1	3	10195	10192	10199	
0	6715	7	1	3	10241	10239	10200	
0	6718	7	1	3	10230	8972	9338	
0	6719	7	1	3	9839	9873	6469	
0	6720	7	1	3	9819	10212	6470	
0	6721	7	1	3	9841	9880	6471	
0	6722	7	1	3	9822	10214	6472	
3	6724	6	0	2	6477	6235	
0	6739	5	1	1	10066	
0	6740	5	1	1	10004	
0	6741	5	1	1	9981	
0	6744	5	1	1	10067	
0	6745	5	1	1	10005	
0	6746	5	1	1	9982	
0	6751	5	1	1	10074	
0	6752	5	1	1	10059	
0	6753	5	1	1	10013	
0	6754	5	1	1	10045	
0	6755	5	1	1	10046	
2	8735	1	523			
0	6760	5	1	1	10075	
0	6761	5	1	1	10060	
0	6762	5	1	1	10014	
0	6772	5	1	1	10177	
0	6773	5	1	1	10130	
0	6776	5	1	1	10178	
0	6777	5	1	1	10131	
0	6782	5	1	1	10170	
0	6783	5	1	1	10139	
0	6784	5	1	1	10156	
0	6785	5	1	1	10157	
0	6790	5	1	1	10171	
0	6791	5	1	1	10140	
0	6792	6	2	2	6630	6631	
0	6795	6	2	2	6632	6633	
0	6801	7	1	2	10222	10247	
0	6802	7	1	2	10252	10226	
0	6803	7	1	2	10243	10218	
0	6804	7	1	2	10232	10256	
0	6805	5	1	1	6466	
0	6806	6	1	2	8135	6651	
0	6807	5	1	1	10263	
0	6808	6	1	2	10264	6653	
0	6809	5	1	1	10265	
0	6810	6	1	2	10266	6655	
0	6811	5	1	1	10267	
0	6812	6	1	2	10268	6657	
0	6813	5	1	1	10269	
0	6814	6	1	2	10270	6659	
0	6815	6	1	2	9824	6661	
0	6816	6	1	2	9672	6663	
0	6817	3	5	2	10244	6664	
2	9497	1	3887			
0	6823	5	1	1	10271	
0	6824	6	1	2	10272	6666	
0	6825	5	1	1	10273	
0	6826	6	1	2	10274	6668	
0	6827	5	1	1	10275	
0	6828	6	1	2	10276	6670	
0	6829	5	1	1	10277	
0	6830	6	1	2	10278	6672	
0	6831	5	2	1	10248	
0	6834	5	1	1	10291	
0	6835	6	1	2	10292	5618	
0	6836	5	1	1	10293	
0	6837	6	1	2	10294	5619	
0	6838	5	1	1	10295	
0	6839	6	1	2	10296	5620	
0	6840	5	1	1	10297	
0	6841	6	1	2	10298	5621	
0	6842	6	1	2	9830	6690	
0	6843	6	1	2	9753	6692	
0	6844	3	5	2	10253	6693	
0	6850	5	1	1	10299	
0	6851	6	1	2	10300	6695	
0	6852	5	1	1	10301	
0	6853	6	1	2	10302	6434	
0	6854	5	1	1	10303	
0	6855	6	1	2	10304	6698	
0	6856	6	1	2	9886	6700	
0	6857	5	2	1	10257	
0	6860	7	1	3	10236	10186	6708	
0	6861	7	1	3	10183	10238	6709	
0	6862	7	1	3	10240	10196	6710	
0	6863	7	1	3	10193	10242	6711	
0	6866	3	5	3	4197	6718	3785	
0	6872	4	1	2	6719	6473	
0	6873	4	1	2	6720	6474	
0	6874	4	1	2	6721	6475	
0	6875	4	1	2	6722	6476	
0	6876	5	1	1	10319	
0	6879	7	1	2	10216	10261	
0	6880	7	1	2	10262	8201	
0	6881	3	2	2	10245	6137	
0	6884	5	1	1	10279	
0	6885	5	2	1	10246	
0	6888	5	1	1	10281	
0	6889	5	1	1	10283	
0	6890	6	1	2	10284	5176	
0	6891	3	2	2	10250	6138	
0	6894	5	1	1	10285	
0	6895	5	1	1	10287	
0	6896	6	1	2	10288	5728	
0	6897	5	2	1	10251	
2	8209	1	137			
0	6900	5	1	1	10289	
0	6901	3	2	2	10254	6193	
0	6904	5	1	1	10305	
0	6905	5	2	1	10255	
0	6908	5	1	1	10307	
0	6909	3	2	2	10259	6194	
0	6912	5	1	1	10309	
0	6913	5	1	1	10311	
0	6914	5	1	1	10313	
0	6915	6	1	2	10314	5734	
0	6916	5	2	1	10260	
0	6919	5	1	1	10315	
0	6922	5	1	1	10317	
0	6923	6	1	2	10318	6067	
3	6924	3	0	2	6382	6801	
3	6925	3	0	2	6386	6802	
3	6926	3	0	2	6388	6803	
3	6927	3	0	2	6392	6804	
0	6930	5	1	1	6724	
0	6932	6	2	2	6650	6806	
0	6935	6	1	2	9901	6807	
0	6936	6	1	2	9902	6809	
0	6937	6	1	2	9913	6811	
2	9520	1	3921			
0	6938	6	1	2	9914	6813	
0	6939	6	1	2	6660	6815	
0	6940	6	1	2	6662	6816	
2	9521	1	3921			
0	6946	6	1	2	9938	6823	
0	6947	6	1	2	9948	6825	
2	9522	1	3921			
0	6948	6	1	2	9959	6827	
0	6949	6	1	2	9969	6829	
2	9523	1	3921			
0	6953	6	1	2	9728	6834	
0	6954	6	1	2	9729	6836	
0	6955	6	1	2	9740	6838	
0	6956	6	1	2	9741	6840	
0	6957	6	1	2	6689	6842	
0	6958	6	1	2	6691	6843	
2	9524	1	3921			
0	6964	6	1	2	10101	6850	
0	6965	6	1	2	9855	6852	
0	6966	6	1	2	10112	6854	
0	6967	6	2	2	6699	6856	
0	6973	4	1	2	6860	6712	
0	6974	4	1	2	6861	6713	
0	6975	4	1	2	6862	6714	
0	6976	4	1	2	6863	6715	
0	6977	5	1	1	10321	
0	6978	5	1	1	10323	
0	6979	3	3	2	6879	6880	
0	6987	6	1	2	9828	6889	
0	6990	6	1	2	9721	6895	
0	6999	6	1	2	9524	6914	
0	7002	6	1	2	9890	6922	
0	7003	6	2	2	6873	6872	
0	7006	6	2	2	6875	6874	
0	7011	7	1	3	10339	9122	9127	
0	7012	7	1	3	10340	9162	9167	
0	7013	7	1	3	10341	9182	9187	
3	7015	5	0	1	10342	
0	7016	7	1	3	10343	9202	9207	
0	7018	6	1	2	6935	6808	
0	7019	6	1	2	6936	6810	
0	7020	6	1	2	6937	6812	
0	7021	6	1	2	6938	6814	
0	7022	5	1	1	6939	
0	7023	5	4	1	10325	
2	8217	1	137			
0	7028	6	2	2	6946	6824	
0	7031	6	2	2	6947	6826	
0	7034	6	2	2	6948	6828	
0	7037	6	2	2	6949	6830	
0	7040	7	1	2	10326	6079	
0	7041	7	2	2	10330	6675	
0	7044	6	1	2	6953	6835	
0	7045	6	1	2	6954	6837	
0	7046	6	1	2	6955	6839	
0	7047	6	1	2	6956	6841	
0	7048	5	1	1	6957	
0	7049	5	4	1	10332	
0	7054	6	2	2	6964	6851	
0	7057	6	2	2	6965	6853	
0	7060	6	2	2	6966	6855	
0	7064	7	1	2	10333	6139	
0	7065	7	2	2	10337	6703	
0	7072	5	1	1	10344	
0	7073	6	1	2	10345	5172	
0	7074	5	1	1	10346	
0	7075	6	1	2	10347	5727	
0	7076	6	2	2	6890	6987	
0	7079	5	1	1	10348	
0	7080	6	2	2	6896	6990	
0	7083	5	1	1	10350	
0	7084	5	1	1	10352	
0	7085	6	1	2	10353	5198	
0	7086	5	1	1	10354	
0	7087	6	1	2	10355	5731	
0	7088	5	1	1	10356	
0	7089	6	1	2	10357	6912	
0	7090	6	2	2	6915	6999	
0	7093	5	1	1	10358	
0	7094	6	2	2	6974	6973	
0	7097	6	2	2	6976	6975	
0	7101	6	2	2	7002	6923	
0	7105	5	1	1	10360	
0	7110	5	1	1	10362	
0	7114	7	1	3	10364	8875	9094	
0	7115	5	1	1	7019	
0	7116	5	1	1	7021	
0	7125	7	1	2	10327	7018	
0	7126	7	1	2	10328	7020	
0	7127	7	1	2	10329	7022	
0	7130	5	1	1	7045	
2	8664	1	457			
0	7131	5	1	1	7047	
0	7139	7	1	2	10334	7044	
0	7140	7	1	2	10335	7046	
0	7141	7	1	2	10336	7048	
0	7146	7	1	3	10361	8973	9318	
0	7147	7	1	3	10363	8974	9339	
0	7149	5	1	1	10367	
0	7150	5	1	1	10369	
0	7151	6	1	2	10370	6876	
0	7152	6	1	2	9826	7072	
0	7153	6	1	2	9699	7074	
0	7158	6	1	2	9832	7084	
0	7159	6	1	2	9797	7086	
0	7160	6	1	2	10310	7088	
0	7166	5	1	1	10381	
0	7167	5	1	1	10379	
0	7168	5	1	1	10377	
0	7169	5	1	1	10375	
0	7170	5	1	1	10393	
0	7171	5	1	1	10391	
0	7172	5	1	1	10389	
0	7173	7	1	2	7115	10371	
0	7174	7	1	2	7116	10372	
0	7175	7	1	2	6940	10373	
0	7176	7	1	2	9931	10374	
0	7177	5	1	1	10383	
0	7178	7	1	2	7130	10385	
0	7179	7	1	2	7131	10386	
0	7180	7	1	2	6958	10387	
0	7181	7	1	2	10094	10388	
0	7182	5	1	1	10395	
0	7183	5	1	1	10403	
0	7184	6	1	2	10404	6977	
0	7185	5	1	1	10405	
0	7186	6	1	2	10406	6978	
0	7187	7	1	3	10382	8975	9319	
0	7188	7	1	3	10380	8976	9320	
0	7189	7	1	3	10378	8977	9321	
0	7190	3	5	3	4956	7146	3781	
0	7196	7	1	3	10394	8978	9340	
0	7197	7	1	3	10392	8979	9341	
0	7198	3	5	3	4960	7147	3786	
0	7204	6	1	2	10407	7149	
0	7205	5	1	1	10408	
0	7206	6	1	2	10320	7150	
0	7207	7	1	3	10376	8980	9359	
0	7208	7	1	3	10390	8981	9379	
0	7209	6	2	2	7073	7152	
0	7212	6	2	2	7075	7153	
2	9575	1	3962			
0	7215	5	1	1	10397	
0	7216	6	1	2	10398	7079	
0	7217	5	1	1	10399	
0	7218	6	1	2	10400	7083	
2	9576	1	3962			
0	7219	6	2	2	7085	7158	
0	7222	6	2	2	7087	7159	
0	7225	6	2	2	7089	7160	
0	7228	5	1	1	10401	
0	7229	6	1	2	10402	7093	
0	7236	3	2	2	7173	7125	
0	7239	3	2	2	7174	7126	
0	7242	3	2	2	7175	7127	
0	7245	3	2	2	7176	7040	
0	7250	3	6	2	7178	7139	
0	7257	3	2	2	7179	7140	
0	7260	3	2	2	7180	7141	
0	7263	3	2	2	7181	7064	
0	7268	6	1	2	10322	7183	
0	7269	6	1	2	10324	7185	
0	7270	3	5	3	4957	7187	3782	
0	7276	3	5	3	4958	7188	3783	
0	7282	3	5	3	4959	7189	3784	
0	7288	3	5	3	4961	7196	3787	
0	7294	3	5	3	3998	7197	3788	
0	7300	6	1	2	10368	7205	
0	7301	6	2	2	7206	7151	
0	7304	3	5	3	4980	7207	3800	
0	7310	3	5	3	4984	7208	3805	
0	7320	6	1	2	10349	7215	
0	7321	6	1	2	10351	7217	
0	7328	6	1	2	10359	7228	
0	7338	7	1	3	10409	8781	9128	
0	7339	7	1	3	10414	9123	9129	
0	7340	7	1	3	10410	8825	9168	
0	7341	7	1	3	10415	9163	9169	
0	7342	7	1	3	10411	8911	9188	
0	7349	7	1	3	10416	9183	9189	
2	10061	1	5536			
0	7357	7	1	3	10417	9203	9208	
3	7363	5	0	1	10418	
0	7364	7	1	3	10412	8933	9209	
3	7365	5	0	1	10413	
2	10062	1	5536			
3	7394	6	0	2	7268	7184	
3	7397	6	0	2	7269	7186	
0	7402	6	2	2	7204	7300	
0	7405	5	1	1	10419	
0	7406	6	1	2	10420	6884	
0	7407	5	1	1	10421	
0	7408	6	1	2	10422	6888	
0	7409	6	2	2	7320	7216	
0	7412	6	2	2	7321	7218	
0	7415	5	1	1	10423	
0	7416	6	1	2	10424	6904	
0	7417	5	1	1	10425	
0	7418	6	1	2	10426	6908	
0	7419	5	1	1	10427	
0	7420	6	1	2	10428	6913	
0	7421	6	2	2	7328	7229	
0	7424	5	1	1	10435	
0	7425	5	1	1	10433	
2	9617	1	4147			
0	7426	5	1	1	10431	
0	7427	5	1	1	10429	
0	7428	5	1	1	10447	
0	7429	5	1	1	10445	
0	7430	5	1	1	10443	
3	7432	5	0	1	10438	
0	7431	5	1	1	10437	
0	7433	7	1	3	10481	9102	9107	
0	7434	7	1	3	10476	8782	9108	
0	7435	3	1	4	7011	7338	3621	2591	
0	7436	7	1	3	10449	8783	9130	
0	7437	7	1	3	10464	9124	9131	
0	7438	7	1	3	10454	8784	9132	
0	7439	7	1	3	10469	9125	9133	
0	7440	7	1	3	10459	8785	9134	
0	7441	7	1	3	10482	9142	9147	
0	7442	7	1	3	10477	8826	9148	
0	7443	3	1	4	7012	7340	3632	2600	
0	7444	7	1	3	10450	8827	9170	
0	7445	7	1	3	10465	9164	9171	
0	7446	7	1	3	10455	8828	9172	
0	7447	7	1	3	10470	9165	9173	
3	7449	3	0	4	7013	7342	3641	2605	
0	7448	7	1	3	10460	8829	9174	
0	7450	7	1	3	10483	9263	9268	
0	7451	7	1	3	10478	8912	9269	
0	7452	7	1	3	10471	9184	9190	
0	7453	7	1	3	10461	8913	9191	
0	7454	7	1	3	10466	9185	9192	
0	7455	7	1	3	10456	8914	9193	
0	7456	7	1	3	10451	8915	9194	
0	7457	7	1	3	10484	9289	9294	
0	7458	7	1	3	10479	8934	9295	
0	7459	7	1	3	10472	9204	9210	
0	7460	7	1	3	10462	8935	9211	
0	7461	7	1	3	10467	9205	9212	
0	7462	7	1	3	10457	8936	9213	
0	7463	7	1	3	10452	8937	9214	
3	7465	5	0	1	10485	
3	7466	5	0	1	10473	
3	7467	5	0	1	10468	
0	7464	7	1	3	10439	8876	8873	
3	7469	3	0	4	7016	7364	3660	2626	
3	7470	5	0	1	10480	
3	7471	5	0	1	10463	
3	7472	5	0	1	10458	
3	7473	5	0	1	10453	
0	7468	5	1	1	10474	
0	7479	7	1	2	10475	9282	
0	7481	7	1	3	10436	8982	9360	
0	7482	7	1	3	10434	8983	9361	
0	7483	7	1	3	10432	8984	9362	
0	7484	7	1	3	10430	8985	9363	
0	7485	7	1	3	10448	8986	9380	
2	9629	1	4200			
0	7486	7	1	3	10446	8987	9381	
0	7487	7	1	3	10444	8988	9382	
0	7488	7	1	3	10440	8989	9383	
0	7489	6	2	2	10365	10441	
0	7492	6	1	2	10280	7405	
0	7493	6	1	2	10282	7407	
2	9631	1	4203			
0	7498	6	1	2	10306	7415	
0	7499	6	1	2	10308	7417	
0	7500	6	1	2	10312	7419	
3	7503	7	0	9	7105	7166	7167	7168	7169	7424	7425	7426	7427	
3	7504	7	0	9	6640	7110	7170	7171	7172	7428	7429	7430	7431	
0	7505	3	1	4	7433	7434	3616	2585	
3	7506	7	0	2	7435	8202	
0	7507	3	1	4	7339	7436	3622	2592	
0	7508	3	1	4	7437	7438	3623	2593	
0	7509	3	1	4	7439	7440	3624	2594	
0	7510	3	1	4	7441	7442	3627	2595	
3	7511	7	0	2	7443	8203	
0	7512	3	1	4	7341	7444	3633	2601	
0	7513	3	1	4	7445	7446	3634	2602	
0	7514	3	1	4	7447	7448	3635	2603	
3	7515	3	0	4	7450	7451	3646	2610	
3	7516	3	0	4	7452	7453	3647	2611	
3	7517	3	0	4	7454	7455	3648	2612	
3	7518	3	0	4	7349	7456	3649	2613	
3	7519	3	0	4	7457	7458	3654	2618	
3	7520	3	0	4	7459	7460	3655	2619	
3	7521	3	0	4	7461	7462	3656	2620	
3	7522	3	0	4	7357	7463	3657	2621	
0	7525	3	1	4	4741	7114	2624	7464	
0	7526	7	1	3	7468	9333	9342	
0	7527	5	1	1	7394	
0	7528	5	1	1	7397	
0	7529	5	1	1	10486	
0	7530	7	1	2	10487	9283	
0	7531	3	5	3	4981	7481	3801	
0	7537	3	5	3	4982	7482	3802	
0	7543	3	5	3	4983	7483	3803	
0	7549	3	5	3	5165	7484	3804	
0	7555	3	5	3	4985	7485	3806	
0	7561	3	5	3	4986	7486	3807	
2	9645	1	4243			
0	7567	3	5	3	4547	7487	3808	
0	7573	3	5	3	4987	7488	3809	
0	7579	6	2	2	7492	7406	
0	7582	6	2	2	7493	7408	
0	7585	5	1	1	10488	
0	7586	6	1	2	10489	6894	
0	7587	5	1	1	10490	
0	7588	6	1	2	10491	6900	
0	7589	6	2	2	7498	7416	
0	7592	6	2	2	7499	7418	
0	7595	6	2	2	7500	7420	
0	7598	5	1	1	10492	
0	7599	6	1	2	10493	6919	
3	7600	7	0	2	7505	8204	
3	7601	7	0	2	7507	8205	
3	7602	7	0	2	7508	8206	
3	7603	7	0	2	7509	8207	
3	7604	7	0	2	7510	8208	
3	7605	7	0	2	7512	8209	
3	7606	7	0	2	7513	8210	
3	7607	7	0	2	7514	8211	
0	7624	7	1	2	10366	10494	
0	7625	7	1	2	10495	10442	
3	7626	7	0	2	1149	7525	
0	7631	7	1	5	8764	7527	7528	6805	6930	
0	7636	7	1	3	7529	9313	9322	
0	7657	6	1	2	10286	7585	
0	7658	6	1	2	10290	7587	
0	7665	6	1	2	10316	7598	
0	7666	7	1	3	10516	9103	9109	
0	7667	7	1	3	10496	8786	9110	
0	7668	7	1	3	10521	9104	9111	
0	7669	7	1	3	10501	8787	9112	
0	7670	7	1	3	10526	9105	9113	
0	7671	7	1	3	10506	8788	9114	
0	7672	7	1	3	10531	9106	9115	
0	7673	7	1	3	10511	8789	9116	
0	7674	7	1	3	10517	9143	9149	
0	7675	7	1	3	10497	8830	9150	
0	7676	7	1	3	10522	9144	9151	
0	7677	7	1	3	10502	8831	9152	
0	7678	7	1	3	10527	9145	9153	
0	7679	7	1	3	10507	8832	9154	
0	7680	7	1	3	10532	9146	9155	
0	7681	7	1	3	10512	8833	9156	
0	7682	7	1	3	10533	9290	9296	
0	7683	7	1	3	10513	8938	9297	
0	7684	7	1	3	10534	9264	9270	
0	7685	7	1	3	10514	8916	9271	
0	7686	7	1	3	10528	9265	9272	
0	7687	7	1	3	10508	8917	9273	
0	7688	7	1	3	10523	9266	9274	
0	7689	7	1	3	10503	8918	9275	
0	7690	7	1	3	10518	9267	9276	
0	7691	7	1	3	10498	8919	9277	
0	7692	7	1	3	10529	9291	9298	
0	7693	7	1	3	10509	8939	9299	
0	7694	7	1	3	10524	9292	9300	
0	7695	7	1	3	10504	8940	9301	
0	7696	7	1	3	10519	9293	9302	
0	7697	7	1	3	10499	8941	9303	
3	7698	3	0	2	7624	7625	
3	7699	5	0	1	10535	
3	7700	5	0	1	10530	
3	7701	5	0	1	10525	
3	7702	5	0	1	10520	
3	7703	7	0	3	1156	7631	8343	
3	7704	5	0	1	10515	
3	7705	5	0	1	10510	
3	7706	5	0	1	10505	
3	7707	5	0	1	10500	
2	9672	1	4290			
0	7708	5	1	1	10536	
0	7709	6	1	2	10537	6739	
0	7710	5	1	1	10538	
0	7711	6	1	2	10539	6744	
0	7712	6	2	2	7657	7586	
0	7715	6	2	2	7658	7588	
0	7718	5	1	1	10540	
0	7719	6	1	2	10541	6772	
0	7720	5	1	1	10542	
0	7721	6	1	2	10543	6776	
0	7722	5	1	1	10544	
0	7723	6	1	2	10545	5733	
0	7724	6	2	2	7665	7599	
0	7727	3	1	4	7666	7667	3617	2586	
2	9677	1	4301			
0	7728	3	1	4	7668	7669	3618	2587	
0	7729	3	1	4	7670	7671	3619	2588	
0	7730	3	1	4	7672	7673	3620	2589	
0	7731	3	1	4	7674	7675	3628	2596	
0	7732	3	1	4	7676	7677	3629	2597	
0	7733	3	1	4	7678	7679	3630	2598	
3	7735	3	0	4	7682	7683	3638	2604	
3	7736	3	0	4	7684	7685	3642	2606	
3	7737	3	0	4	7686	7687	3643	2607	
3	7738	3	0	4	7688	7689	3644	2608	
3	7739	3	0	4	7690	7691	3645	2609	
3	7740	3	0	4	7692	7693	3651	2615	
3	7741	3	0	4	7694	7695	3652	2616	
3	7742	3	0	4	7696	7697	3653	2617	
0	7734	3	1	4	7680	7681	3631	2599	
0	7743	6	1	2	10068	7708	
0	7744	6	1	2	10069	7710	
2	9195	1	2790			
0	7749	6	1	2	10179	7718	
0	7750	6	1	2	10180	7720	
0	7751	6	1	2	9815	7722	
3	7754	7	0	2	7727	8212	
3	7755	7	0	2	7728	8213	
3	7756	7	0	2	7729	8214	
3	7757	7	0	2	7730	8215	
3	7758	7	0	2	7731	8216	
3	7759	7	0	2	7732	8217	
3	7760	7	0	2	7733	8218	
3	7761	7	0	2	7734	8219	
0	7762	6	2	2	7743	7709	
0	7765	6	2	2	7744	7711	
0	7768	5	1	1	10546	
0	7769	6	1	2	10547	6751	
0	7770	5	1	1	10548	
0	7771	6	1	2	10549	6760	
0	7772	6	2	2	7749	7719	
0	7775	6	2	2	7750	7721	
0	7778	6	2	2	7751	7723	
0	7781	5	1	1	10550	
0	7782	6	1	2	10551	5735	
2	9688	1	4316			
0	7787	6	1	2	10076	7768	
2	9689	1	4316			
0	7788	6	1	2	10077	7770	
0	7795	6	1	2	9816	7781	
0	7796	5	1	1	10552	
0	7797	6	1	2	10553	6740	
0	7798	5	1	1	10554	
0	7799	6	1	2	10555	6745	
0	7800	6	2	2	7787	7769	
0	7803	6	2	2	7788	7771	
0	7806	5	1	1	10556	
0	7807	6	1	2	10557	6773	
0	7808	5	1	1	10558	
0	7809	6	1	2	10559	6777	
0	7810	5	1	1	10560	
0	7811	6	1	2	10561	6782	
0	7812	6	2	2	7795	7782	
0	7815	6	1	2	10006	7796	
0	7816	6	1	2	10007	7798	
0	8126	7	1	2	8122	8221	
0	7821	6	1	2	10132	7806	
0	7822	6	1	2	10133	7808	
0	7823	6	1	2	10172	7810	
0	7826	6	2	2	7815	7797	
0	7829	6	2	2	7816	7799	
0	7832	5	1	1	10562	
0	7833	6	1	2	10563	6752	
0	7834	5	1	1	10564	
0	7835	6	1	2	10565	6761	
0	7836	6	2	2	7821	7807	
0	7839	6	2	2	7822	7809	
0	7842	6	2	2	7823	7811	
0	7845	5	1	1	10566	
0	7846	6	1	2	10567	6790	
0	7851	6	1	2	10061	7832	
0	7852	6	1	2	10062	7834	
0	7859	6	1	2	10173	7845	
0	7860	5	1	1	10568	
0	7861	6	1	2	10569	6741	
0	7862	5	1	1	10570	
0	7863	6	1	2	10571	6746	
0	7864	6	2	2	7851	7833	
0	7867	6	2	2	7852	7835	
0	7870	5	1	1	10572	
0	7871	6	1	2	10573	5730	
0	7872	5	1	1	10574	
0	7873	6	1	2	10575	5732	
0	7874	5	1	1	10576	
0	7875	6	1	2	10577	6783	
0	7876	6	2	2	7859	7846	
0	7879	6	1	2	9983	7860	
0	7880	6	1	2	9984	7862	
0	7885	6	1	2	9774	7870	
0	7886	6	1	2	9775	7872	
0	7887	6	1	2	10141	7874	
0	7890	6	2	2	7879	7861	
0	7893	6	2	2	7880	7863	
0	7896	5	1	1	10578	
0	7897	6	1	2	10579	6753	
0	7898	5	1	1	10580	
0	7899	6	1	2	10581	6762	
0	7900	6	2	2	7885	7871	
0	7903	6	2	2	7886	7873	
0	7906	6	2	2	7887	7875	
0	7909	5	1	1	10582	
0	7910	6	1	2	10583	6791	
0	7917	6	1	2	10015	7896	
0	7918	6	1	2	10016	7898	
0	7923	6	1	2	10142	7909	
0	7924	5	1	1	10584	
0	7925	6	1	2	10585	6680	
0	7926	5	1	1	10586	
0	7927	6	1	2	10587	6681	
0	7928	5	1	1	10588	
0	7929	6	1	2	10589	5690	
0	7930	5	1	1	10590	
0	7931	6	1	2	10591	5691	
0	7932	6	2	2	7917	7897	
0	7935	6	2	2	7918	7899	
0	7938	5	1	1	10592	
0	7939	6	1	2	10593	6784	
0	7940	6	2	2	7923	7910	
0	7943	6	1	2	9995	7924	
0	7944	6	1	2	9996	7926	
0	7945	6	1	2	9786	7928	
0	7946	6	1	2	9787	7930	
0	7951	6	1	2	10158	7938	
0	7954	6	2	2	7943	7925	
0	7957	6	2	2	7944	7927	
0	7960	6	2	2	7945	7929	
0	7963	6	2	2	7946	7931	
0	7966	5	1	1	10594	
0	7967	6	1	2	10595	6754	
0	7968	5	1	1	10596	
0	7969	6	1	2	10597	6755	
0	7970	6	2	2	7951	7939	
2	9760	1	4400			
0	7973	5	1	1	10598	
0	7974	6	1	2	10599	6785	
0	7984	6	1	2	10047	7966	
0	7985	6	1	2	10048	7968	
0	7987	6	1	2	10159	7973	
0	7988	7	1	3	10602	10331	9071	
0	7989	7	1	3	10600	10249	9072	
0	7990	7	1	3	10603	10384	8766	
2	10158	1	5655			
0	7991	7	1	3	10601	7177	8767	
0	7992	5	1	1	10608	
0	7993	6	1	2	10609	6448	
0	7994	7	1	3	10606	10338	9074	
0	7995	7	1	3	10604	10258	9075	
0	7996	7	1	3	10607	10396	8858	
0	7997	7	1	3	10605	7182	8859	
0	7998	6	2	2	7984	7967	
0	8001	6	2	2	7985	7969	
0	8004	6	2	2	7987	7974	
0	8009	6	1	2	9869	7992	
0	8013	3	2	4	7988	7989	7990	7991	
0	8017	3	2	4	7994	7995	7996	7997	
0	8020	5	1	1	10610	
0	8021	6	1	2	10611	6682	
0	8022	5	1	1	10612	
0	8023	6	1	2	10613	6683	
0	8025	6	1	2	8009	7993	
0	8026	5	1	1	10614	
0	8027	6	1	2	10615	6449	
0	8031	6	1	2	10030	8020	
0	8032	6	1	2	10031	8022	
0	8033	5	1	1	10616	
0	8034	6	1	2	9870	8026	
0	8035	7	1	2	8860	8025	
0	8036	5	1	1	10618	
0	8037	6	1	2	8031	8021	
0	8038	6	1	2	8032	8023	
0	8039	6	1	2	8034	8027	
0	8040	5	1	1	8038	
0	8041	7	1	2	8768	8037	
0	8042	5	1	1	8039	
0	8043	7	1	2	8040	9073	
0	8044	7	1	2	8042	9076	
0	8045	3	2	2	8043	8041	
0	8048	3	2	2	8044	8035	
2	9741	1	4364			
0	8055	6	1	2	10620	8033	
0	8056	5	1	1	10621	
0	8057	6	1	2	10622	8036	
0	8058	5	1	1	10623	
0	8059	6	1	2	10617	8056	
0	8060	6	1	2	10619	8058	
0	8061	6	2	2	8055	8059	
0	8064	6	2	2	8057	8060	
0	8071	7	1	3	10626	8990	9343	
0	8072	7	1	3	10624	8991	9323	
0	8073	5	1	1	10625	
0	8074	5	1	1	10627	
3	8075	3	0	4	7526	8071	3659	2625	
3	8076	3	0	4	7636	8072	3661	2627	
2	9746	1	4379			
0	8077	7	1	2	8073	8992	
0	8078	7	1	2	8074	8993	
0	8079	3	2	2	7530	8077	
0	8082	3	2	2	7479	8078	
0	8089	7	1	2	10628	9278	
0	8090	7	1	2	10630	9279	
0	8091	7	1	2	10629	9280	
0	8092	7	1	2	10631	9281	
0	8093	3	2	2	8089	3071	
0	8096	3	2	2	8090	3072	
0	8099	3	2	2	8091	3073	
0	8102	3	2	2	8092	3074	
2	9753	1	4385			
0	8113	7	1	3	10638	9186	9195	
0	8114	7	1	3	10636	8920	9196	
0	8115	7	1	3	10639	9206	9215	
2	10159	1	5655			
0	8116	7	1	3	10637	8942	9216	
0	8117	7	1	3	10634	9126	9135	
0	8118	7	1	3	10632	8790	9136	
0	8119	7	1	3	10635	9166	9175	
0	8120	7	1	3	10633	8834	9176	
0	8121	3	1	4	8117	8118	3662	2703	
3	8123	3	0	4	8113	8114	3650	2614	
3	8124	3	0	4	8115	8116	3658	2622	
0	8122	3	1	4	8119	8120	3663	2778	
0	8125	7	1	2	8121	8220	
3	8127	5	0	1	8125	
3	8128	5	0	1	8126	
2	8129	1	4			
2	8130	1	4			
2	8131	1	4			
2	8132	1	4			
2	8133	1	4			
2	8134	1	4			
2	8135	1	4			
2	8136	1	11			
2	8137	1	11			
2	8138	1	14			
2	8139	1	14			
2	8140	1	17			
2	8141	1	17			
2	8142	1	20			
2	8143	1	20			
2	8144	1	27			
2	8145	1	27			
2	8146	1	27			
2	8147	1	31			
2	8148	1	31			
2	8149	1	34			
2	8150	1	34			
2	8151	1	37			
2	8152	1	37			
2	8153	1	40			
2	8154	1	40			
2	8155	1	43			
2	8156	1	43			
2	8157	1	46			
2	8158	1	46			
2	8159	1	49			
2	8160	1	49			
2	8161	1	54			
2	8162	1	54			
2	8163	1	54			
2	8164	1	54			
2	8165	1	54			
2	8166	1	54			
2	8167	1	54			
2	8168	1	61			
2	8169	1	61			
2	8170	1	64			
2	8171	1	64			
2	8172	1	67			
2	8173	1	67			
2	8174	1	70			
2	8175	1	70			
2	8176	1	73			
2	8177	1	73			
2	8178	1	76			
2	8179	1	76			
2	8180	1	83			
2	8181	1	83			
2	8182	1	88			
2	8183	1	88			
2	8184	1	91			
2	8185	1	91			
2	8186	1	94			
2	8187	1	94			
2	8188	1	97			
2	8189	1	97			
2	8190	1	100			
2	8191	1	100			
