1 N1 0 2 0
1 N4 0 3 0
1 N8 0 3 0
1 N11 0 2 0
1 N14 0 2 0
1 N17 0 3 0
1 N21 0 1 0
1 N24 0 1 0
1 N27 0 2 0
1 N30 0 2 0
1 N34 0 2 0
1 N37 0 2 0
1 N40 0 2 0
1 N43 0 2 0
1 N47 0 2 0
1 N50 0 2 0
1 N53 0 2 0
1 N56 0 2 0
1 N60 0 1 0
1 N63 0 2 0
1 N66 0 2 0
1 N69 0 2 0
1 N73 0 1 0
1 N76 0 2 0
1 N79 0 2 0
1 N82 0 2 0
1 N86 0 2 0
1 N89 0 2 0
1 N92 0 1 0
1 N95 0 2 0
1 N99 0 1 0
1 N102 0 2 0
1 N105 0 1 0
1 N108 0 3 0
1 N112 0 1 0
1 N115 0 1 0
0 n214 5 2 1 N92
0 n206 5 2 1 N105
0 n208 5 2 1 N99
0 n226 5 2 1 N21
0 n219 5 2 1 N73
0 n231 5 2 1 N60
2 N1-1 1 N1 
2 N1-2 1 N1 
2 N4-1 1 N4 
2 N4-2 1 N4 
2 N4-3 1 N4 
2 N8-1 1 N8 
2 N8-2 1 N8 
2 N8-3 1 N8 
2 N11-1 1 N11 
2 N11-2 1 N11 
2 N14-1 1 N14 
2 N14-2 1 N14 
2 N17-1 1 N17 
2 N17-2 1 N17 
2 N17-3 1 N17 
2 N27-1 1 N27 
2 N27-2 1 N27 
2 N30-1 1 N30 
2 N30-2 1 N30 
2 N34-1 1 N34 
2 N34-2 1 N34 
2 N37-1 1 N37 
2 N37-2 1 N37 
2 N40-1 1 N40 
2 N40-2 1 N40 
2 N43-1 1 N43 
2 N43-2 1 N43 
2 N47-1 1 N47 
2 N47-2 1 N47 
2 N50-1 1 N50 
2 N50-2 1 N50 
2 N53-1 1 N53 
2 N53-2 1 N53 
2 N56-1 1 N56 
2 N56-2 1 N56 
2 N63-1 1 N63 
2 N63-2 1 N63 
2 N66-1 1 N66 
2 N66-2 1 N66 
2 N69-1 1 N69 
2 N69-2 1 N69 
2 N76-1 1 N76 
2 N76-2 1 N76 
2 N79-1 1 N79 
2 N79-2 1 N79 
2 N82-1 1 N82 
2 N82-2 1 N82 
2 N86-1 1 N86 
2 N86-2 1 N86 
2 N89-1 1 N89 
2 N89-2 1 N89 
2 N95-1 1 N95 
2 N95-2 1 N95 
2 N102-1 1 N102 
2 N102-2 1 N102 
2 N108-1 1 N108 
2 N108-2 1 N108 
2 N108-3 1 N108 
0 n235 5 1 1 N53-1
0 n285 5 1 1 N17-1
0 n287 5 2 1 N11-2
0 n326 5 1 1 N37-2
0 n329 5 1 1 N102-2
0 n266 5 2 1 N4-3
0 n241 5 3 1 N30-2
0 n335 5 1 1 N76-2
0 n336 5 1 1 N89-2
0 n339 5 1 1 N50-2
0 n340 5 1 1 N63-2
2 n214-1 1 n214 
2 n214-2 1 n214 
2 n206-1 1 n206 
2 n206-2 1 n206 
2 n208-1 1 n208 
2 n208-2 1 n208 
2 n226-1 1 n226 
2 n226-2 1 n226 
2 n219-1 1 n219 
2 n219-2 1 n219 
2 n231-1 1 n231 
2 n231-2 1 n231 
0 n324 6 1 2 n326 N43-2
0 n328 6 1 2 n329 N108-3
0 n334 6 1 2 n335 N82-2
0 n333 6 1 2 n336 N95-2
0 n338 6 1 2 n339 N56-2
0 n337 6 1 2 n340 N69-2
2 n287-1 1 n287 
2 n287-2 1 n287 
2 n266-1 1 n266 
2 n266-2 1 n266 
2 n241-1 1 n241 
2 n241-2 1 n241 
2 n241-3 1 n241 
0 n325 6 1 2 N17-3 n287-2
0 n330 4 1 2 N1-2 n266-2
0 n318 4 2 2 N24 n241-3
0 n332 6 1 2 n333 n334
0 n331 6 1 2 n337 n338
0 n323 6 1 2 n324 n325
0 n320 4 1 2 n331 n332
2 n318-1 1 n318 
2 n318-2 1 n318 
0 n327 4 1 2 n330 n318-2
0 n322 6 1 2 n327 n328
0 n321 4 1 2 n322 n323
3 N223 6 0 2 n320 n321
2 N223-1 1 N223 
2 N223-2 1 N223 
2 N223-3 1 N223 
2 N223-4 1 N223 
2 N223-5 1 N223 
2 N223-6 1 N223 
2 N223-7 1 N223 
2 N223-8 1 N223 
2 N223-9 1 N223 
0 n304 6 1 2 N89-1 N223-1
0 n305 6 1 2 N11-1 N223-2
0 n308 6 1 2 N102-1 N223-3
0 n309 6 1 2 N63-1 N223-4
0 n310 6 1 2 N76-1 N223-5
0 n315 6 1 2 N37-1 N223-6
0 n246 6 2 2 N1-1 N223-7
0 n286 5 2 1 N223-8
0 n319 6 1 2 N50-1 N223-9
0 n272 6 2 2 n304 N95-1
0 n223 7 2 2 n305 N17-2
0 n255 6 2 2 n308 N108-2
0 n216 7 3 2 n309 N69-1
0 n211 6 3 2 n310 N82-1
0 n188 6 3 2 n315 N43-1
0 n228 7 3 2 n319 N56-1
2 n246-1 1 n246 
2 n246-2 1 n246 
2 n286-1 1 n286 
2 n286-2 1 n286 
0 n284 4 1 2 n286-1 n287-1
0 n264 5 2 1 n246-2
0 n238 4 3 2 n286-2 n318-1
2 n272-1 1 n272 
2 n272-2 1 n272 
2 n223-1 1 n223 
2 n223-2 1 n223 
2 n255-1 1 n255 
2 n255-2 1 n255 
2 n216-1 1 n216 
2 n216-2 1 n216 
2 n216-3 1 n216 
2 n211-1 1 n211 
2 n211-2 1 n211 
2 n211-3 1 n211 
2 n188-1 1 n188 
2 n188-2 1 n188 
2 n188-3 1 n188 
2 n228-1 1 n228 
2 n228-2 1 n228 
2 n228-3 1 n228 
0 n254 5 1 1 n255-1
0 n233 5 2 1 n188-2
0 n280 4 1 2 n284 n285
0 n202 5 2 1 n272-2
0 n283 6 2 2 n226-2 n223-2
0 n257 4 2 2 N112 n255-2
0 n296 7 2 2 n219-2 n216-3
0 n271 4 2 2 N86-2 n211-3
0 n187 4 3 2 N47-2 n188-3
0 n299 6 2 2 n231-2 n228-3
2 n264-1 1 n264 
2 n264-2 1 n264 
2 n238-1 1 n238 
2 n238-2 1 n238 
2 n238-3 1 n238 
0 n263 4 1 2 N14-2 n264-1
0 n289 4 1 2 N40-2 n238-2
0 n316 4 1 2 N8-3 n264-2
0 n317 4 1 2 N34-2 n238-3
2 n233-1 1 n233 
2 n233-2 1 n233 
2 n202-1 1 n202 
2 n202-2 1 n202 
2 n283-1 1 n283 
2 n283-2 1 n283 
2 n257-1 1 n257 
2 n257-2 1 n257 
2 n296-1 1 n296 
2 n296-2 1 n296 
2 n271-1 1 n271 
2 n271-2 1 n271 
2 n187-1 1 n187 
2 n187-2 1 n187 
2 n187-3 1 n187 
2 n299-1 1 n299 
2 n299-2 1 n299 
0 n275 6 2 2 n208-2 n202-2
0 n307 5 1 1 n257-2
0 n306 4 1 2 n296-2 n271-2
0 n314 5 1 1 n187-3
0 n313 6 1 2 n316 N4-2
0 n291 6 2 2 n317 N30-1
0 n302 6 1 2 n306 n307
0 n312 6 1 2 n313 n314
2 n275-1 1 n275 
2 n275-2 1 n275 
2 n291-1 1 n291 
2 n291-2 1 n291 
0 n303 6 1 2 n275-2 n283-2
0 n311 6 1 2 n291-2 n299-2
0 n301 4 1 2 n302 n303
0 n300 4 1 2 n311 n312
3 N329 6 0 2 n300 n301
2 N329-1 1 N329 
2 N329-2 1 N329 
2 N329-3 1 N329 
2 N329-4 1 N329 
2 N329-5 1 N329 
2 N329-6 1 N329 
2 N329-7 1 N329 
2 N329-8 1 N329 
2 N329-9 1 N329 
2 N329-10 1 N329 
2 N329-11 1 N329 
0 n186 4 1 2 N329-1 n188-1
0 n212 7 1 2 N86-1 N329-2
0 n234 7 1 2 N47-1 N329-3
0 n239 7 1 2 N34-1 N329-4
0 n245 6 1 2 N8-1 N329-5
0 n265 7 1 2 N8-2 N329-6
0 n274 6 1 2 N329-7 n275-1
0 n282 7 1 2 N329-8 n283-1
0 n290 7 1 2 N329-9 n291-1
0 n207 5 8 1 N329-10
0 n298 7 1 2 N329-11 n299-1
0 n184 4 1 2 n186 n187-1
0 n237 4 1 2 n239 n238-1
0 n242 6 1 2 n245 n246-1
0 n262 4 1 2 n265 n266-1
0 n273 6 1 2 n274 n206-2
0 n281 4 1 2 n282 N27-2
0 n288 4 1 2 n290 n241-2
0 n297 4 1 2 n298 N66-2
2 n207-1 1 n207 
2 n207-2 1 n207 
2 n207-3 1 n207 
2 n207-4 1 n207 
2 n207-5 1 n207 
2 n207-6 1 n207 
2 n207-7 1 n207 
2 n207-8 1 n207 
0 n203 4 1 2 n207-1 n208-1
0 n217 4 1 2 n207-2 n219-1
0 n224 4 1 2 n207-3 n226-1
0 n230 4 1 2 n207-4 n231-1
0 n256 4 1 2 n207-5 n257-1
0 n259 4 1 2 n207-6 n187-2
0 n261 6 1 2 n262 n263
0 n270 3 1 2 n207-7 n271-1
0 n267 4 1 2 n273 n272-1
0 n279 6 1 2 n280 n281
0 n278 6 1 2 n288 n289
0 n295 4 1 2 n207-8 n296-1
0 n292 6 1 2 n297 n228-2
0 n253 4 1 2 N115 n256
0 n258 4 1 2 n259 N53-2
0 n269 6 1 2 n270 n214-2
0 n277 6 1 2 n278 n279
0 n294 4 1 2 n295 N79-2
0 n252 6 1 2 n253 n254
0 n251 6 1 2 n258 n233-2
0 n268 4 1 2 n269 n211-2
0 n293 6 1 2 n294 n216-2
0 n250 6 1 2 n251 n252
0 n260 4 1 2 n267 n268
0 n276 6 1 2 n292 n293
0 n249 6 1 2 n260 n261
0 n247 4 1 2 n276 n277
0 n248 4 1 2 n249 n250
3 N370 6 0 2 n247 n248
2 N370-1 1 N370 
2 N370-2 1 N370 
2 N370-3 1 N370 
2 N370-4 1 N370 
2 N370-5 1 N370 
2 N370-6 1 N370 
0 n218 7 1 2 N79-1 N370-1
0 n225 7 1 2 N27-1 N370-2
0 n229 7 1 2 N66-1 N370-3
0 n205 5 3 1 N370-4
0 n240 7 1 2 N40-1 N370-5
0 n244 6 1 2 N14-1 N370-6
0 n215 4 1 2 n217 n218
0 n222 4 1 2 n224 n225
0 n227 4 1 2 n229 n230
0 n236 4 1 2 n240 n241-1
0 n243 6 1 2 n244 N4-1
2 n205-1 1 n205 
2 n205-2 1 n205 
2 n205-3 1 n205 
0 n204 4 1 2 n205-1 n206-1
0 n213 4 1 2 n205-2 n214-1
0 n178 6 2 2 n215 n216-1
0 n172 6 2 2 n222 n223-1
0 n179 7 3 2 n227 n228-1
0 n185 4 2 2 n235 n205-3
0 n175 6 2 2 n236 n237
0 n196 4 1 2 n242 n243
0 n201 4 1 2 n203 n204
0 n210 3 1 2 n212 n213
2 n178-1 1 n178 
2 n178-2 1 n178 
2 n172-1 1 n172 
2 n172-2 1 n172 
2 n179-1 1 n179 
2 n179-2 1 n179 
2 n179-3 1 n179 
2 n185-1 1 n185 
2 n185-2 1 n185 
2 n175-1 1 n175 
2 n175-2 1 n175 
0 n177 3 1 2 n178-1 n179-1
0 n180 4 1 2 n184 n185-1
0 n183 6 2 2 n201 n202-1
0 n182 4 2 2 n210 n211-1
0 n194 5 2 1 n172-2
0 n232 4 1 2 n234 n185-2
0 n195 5 2 1 n175-2
0 n193 7 2 2 n232 n233-1
2 n183-1 1 n183 
2 n183-2 1 n183 
2 n182-1 1 n182 
2 n182-2 1 n182 
2 n194-1 1 n194 
2 n194-2 1 n194 
2 n195-1 1 n195 
2 n195-2 1 n195 
0 n181 4 1 2 n183-1 n182-1
0 n189 4 1 2 n194-1 n195-1
0 n209 5 1 1 n182-2
0 n221 4 1 2 n194-2 n179-3
2 n193-1 1 n193 
2 n193-2 1 n193 
0 n176 4 1 2 n180 n181
0 n191 4 1 2 n179-2 n193-1
0 n192 6 2 2 n209 n178-2
0 n220 4 1 2 n193-2 n195-2
0 n174 6 1 2 n176 n177
3 N430 6 0 2 n220 n221
2 n192-1 1 n192 
2 n192-2 1 n192 
0 n173 6 1 2 n174 n175-1
0 n190 6 1 2 n191 n192-1
0 n200 5 1 1 n192-2
0 n198 3 1 2 N430 N108-1
3 N432 6 0 2 n173 n172-1
3 N431 6 0 2 n189 n190
0 n199 6 1 2 n200 n183-2
0 n197 4 1 2 n198 n199
3 N421 4 0 2 n196 n197
