module c1355(N1,N8,N15,N22,N29,N36,N43,N50,N57,N64,N71,N78,
             N85,N92,N99,N106,N113,N120,N127,N134,N141,N148,
			 N155,N162,N169,N176,N183,N190,N197,N204,N211,N218,
			 N225,N226,N227,N228,N229,N230,N231,N232,N233,N1324,
			 N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,
			 N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
			 N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355);

input N1,N8,N15,N22,N29,N36,N43,N50,N57,N64,N71,N78,N85,N92,N99,N106,N113,N120,N127,N134,
      N141,N148,N155,N162,N169,N176,N183,N190,N197,N204,N211,N218,N225,N226,N227,N228,N229,
	  N230,N231,N232,N233;

output N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,
       N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,
	   N1352,N1353,N1354,N1355;

wire N242,N245,N248,N251,N254,N257,N260,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,
     N293,N296,N299,N302,N305,N308,N311,N314,N317,N320,N323,N326,N329,N332,N335,N338,N341,
	 N344,N347,N350,N353,N356,N359,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
	 N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
	 N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,
	 N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,
	 N424,N425,N426,N429,N432,N435,N438,N441,N444,N447,N450,N453,N456,N459,N462,N465,N468,
	 N471,N474,N477,N480,N483,N486,N489,N492,N495,N498,N501,N504,N507,N510,N513,N516,N519,
	 N522,N525,N528,N531,N534,N537,N540,N543,N546,N549,N552,N555,N558,N561,N564,N567,N570,
	 N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,
	 N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,N612,
	 N617,N622,N627,N632,N637,N642,N645,N648,N651,N654,N657,N660,N663,N666,N669,N672,N675,
	 N678,N681,N684,N687,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
	 N703,N704,N705,N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,N736,N739,N742,N745,
	 N748,N751,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
	 N769,N770,N773,N776,N779,N782,N785,N788,N791,N794,N797,N800,N803,N806,N809,N812,N815,
	 N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
	 N847,N860,N873,N886,N899,N912,N925,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
	 N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,
	 N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
	 N982,N983,N984,N985,N986,N991,N996,N1001,N1006,N1011,N1016,N1021,N1026,N1031,N1036,N1039,
	 N1042,N1045,N1048,N1051,N1054,N1057,N1060,N1063,N1066,N1069,N1072,N1075,N1078,N1081,N1084,
	 N1087,N1090,N1093,N1096,N1099,N1102,N1105,N1108,N1111,N1114,N1117,N1120,N1123,N1126,N1129,
	 N1132,N1135,N1138,N1141,N1144,N1147,N1150,N1153,N1156,N1159,N1162,N1165,N1168,N1171,N1174,
	 N1177,N1180,N1183,N1186,N1189,N1192,N1195,N1198,N1201,N1204,N1207,N1210,N1213,N1216,N1219,
	 N1222,N1225,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,
	 N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,
	 N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,
	 N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
	 N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,
	 N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,
	 N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323;

and AND2_0(N242,N225,N233);
and AND2_1(N245,N226,N233);
and AND2_2(N248,N227,N233);
and AND2_3(N251,N228,N233);
and AND2_4(N254,N229,N233);
and AND2_5(N257,N230,N233);
and AND2_6(N260,N231,N233);
and AND2_7(N263,N232,N233);
nand NAND2_0(N266,N1,N8);
nand NAND2_1(N269,N15,N22);
nand NAND2_2(N272,N29,N36);
nand NAND2_3(N275,N43,N50);
nand NAND2_4(N278,N57,N64);
nand NAND2_5(N281,N71,N78);
nand NAND2_6(N284,N85,N92);
nand NAND2_7(N287,N99,N106);
nand NAND2_8(N290,N113,N120);
nand NAND2_9(N293,N127,N134);
nand NAND2_10(N296,N141,N148);
nand NAND2_11(N299,N155,N162);
nand NAND2_12(N302,N169,N176);
nand NAND2_13(N305,N183,N190);
nand NAND2_14(N308,N197,N204);
nand NAND2_15(N311,N211,N218);
nand NAND2_16(N314,N1,N29);
nand NAND2_17(N317,N57,N85);
nand NAND2_18(N320,N8,N36);
nand NAND2_19(N323,N64,N92);
nand NAND2_20(N326,N15,N43);
nand NAND2_21(N329,N71,N99);
nand NAND2_22(N332,N22,N50);
nand NAND2_23(N335,N78,N106);
nand NAND2_24(N338,N113,N141);
nand NAND2_25(N341,N169,N197);
nand NAND2_26(N344,N120,N148);
nand NAND2_27(N347,N176,N204);
nand NAND2_28(N350,N127,N155);
nand NAND2_29(N353,N183,N211);
nand NAND2_30(N356,N134,N162);
nand NAND2_31(N359,N190,N218);
nand NAND2_32(N362,N1,N266);
nand NAND2_33(N363,N8,N266);
nand NAND2_34(N364,N15,N269);
nand NAND2_35(N365,N22,N269);
nand NAND2_36(N366,N29,N272);
nand NAND2_37(N367,N36,N272);
nand NAND2_38(N368,N43,N275);
nand NAND2_39(N369,N50,N275);
nand NAND2_40(N370,N57,N278);
nand NAND2_41(N371,N64,N278);
nand NAND2_42(N372,N71,N281);
nand NAND2_43(N373,N78,N281);
nand NAND2_44(N374,N85,N284);
nand NAND2_45(N375,N92,N284);
nand NAND2_46(N376,N99,N287);
nand NAND2_47(N377,N106,N287);
nand NAND2_48(N378,N113,N290);
nand NAND2_49(N379,N120,N290);
nand NAND2_50(N380,N127,N293);
nand NAND2_51(N381,N134,N293);
nand NAND2_52(N382,N141,N296);
nand NAND2_53(N383,N148,N296);
nand NAND2_54(N384,N155,N299);
nand NAND2_55(N385,N162,N299);
nand NAND2_56(N386,N169,N302);
nand NAND2_57(N387,N176,N302);
nand NAND2_58(N388,N183,N305);
nand NAND2_59(N389,N190,N305);
nand NAND2_60(N390,N197,N308);
nand NAND2_61(N391,N204,N308);
nand NAND2_62(N392,N211,N311);
nand NAND2_63(N393,N218,N311);
nand NAND2_64(N394,N1,N314);
nand NAND2_65(N395,N29,N314);
nand NAND2_66(N396,N57,N317);
nand NAND2_67(N397,N85,N317);
nand NAND2_68(N398,N8,N320);
nand NAND2_69(N399,N36,N320);
nand NAND2_70(N400,N64,N323);
nand NAND2_71(N401,N92,N323);
nand NAND2_72(N402,N15,N326);
nand NAND2_73(N403,N43,N326);
nand NAND2_74(N404,N71,N329);
nand NAND2_75(N405,N99,N329);
nand NAND2_76(N406,N22,N332);
nand NAND2_77(N407,N50,N332);
nand NAND2_78(N408,N78,N335);
nand NAND2_79(N409,N106,N335);
nand NAND2_80(N410,N113,N338);
nand NAND2_81(N411,N141,N338);
nand NAND2_82(N412,N169,N341);
nand NAND2_83(N413,N197,N341);
nand NAND2_84(N414,N120,N344);
nand NAND2_85(N415,N148,N344);
nand NAND2_86(N416,N176,N347);
nand NAND2_87(N417,N204,N347);
nand NAND2_88(N418,N127,N350);
nand NAND2_89(N419,N155,N350);
nand NAND2_90(N420,N183,N353);
nand NAND2_91(N421,N211,N353);
nand NAND2_92(N422,N134,N356);
nand NAND2_93(N423,N162,N356);
nand NAND2_94(N424,N190,N359);
nand NAND2_95(N425,N218,N359);
nand NAND2_96(N426,N362,N363);
nand NAND2_97(N429,N364,N365);
nand NAND2_98(N432,N366,N367);
nand NAND2_99(N435,N368,N369);
nand NAND2_100(N438,N370,N371);
nand NAND2_101(N441,N372,N373);
nand NAND2_102(N444,N374,N375);
nand NAND2_103(N447,N376,N377);
nand NAND2_104(N450,N378,N379);
nand NAND2_105(N453,N380,N381);
nand NAND2_106(N456,N382,N383);
nand NAND2_107(N459,N384,N385);
nand NAND2_108(N462,N386,N387);
nand NAND2_109(N465,N388,N389);
nand NAND2_110(N468,N390,N391);
nand NAND2_111(N471,N392,N393);
nand NAND2_112(N474,N394,N395);
nand NAND2_113(N477,N396,N397);
nand NAND2_114(N480,N398,N399);
nand NAND2_115(N483,N400,N401);
nand NAND2_116(N486,N402,N403);
nand NAND2_117(N489,N404,N405);
nand NAND2_118(N492,N406,N407);
nand NAND2_119(N495,N408,N409);
nand NAND2_120(N498,N410,N411);
nand NAND2_121(N501,N412,N413);
nand NAND2_122(N504,N414,N415);
nand NAND2_123(N507,N416,N417);
nand NAND2_124(N510,N418,N419);
nand NAND2_125(N513,N420,N421);
nand NAND2_126(N516,N422,N423);
nand NAND2_127(N519,N424,N425);
nand NAND2_128(N522,N426,N429);
nand NAND2_129(N525,N432,N435);
nand NAND2_130(N528,N438,N441);
nand NAND2_131(N531,N444,N447);
nand NAND2_132(N534,N450,N453);
nand NAND2_133(N537,N456,N459);
nand NAND2_134(N540,N462,N465);
nand NAND2_135(N543,N468,N471);
nand NAND2_136(N546,N474,N477);
nand NAND2_137(N549,N480,N483);
nand NAND2_138(N552,N486,N489);
nand NAND2_139(N555,N492,N495);
nand NAND2_140(N558,N498,N501);
nand NAND2_141(N561,N504,N507);
nand NAND2_142(N564,N510,N513);
nand NAND2_143(N567,N516,N519);
nand NAND2_144(N570,N426,N522);
nand NAND2_145(N571,N429,N522);
nand NAND2_146(N572,N432,N525);
nand NAND2_147(N573,N435,N525);
nand NAND2_148(N574,N438,N528);
nand NAND2_149(N575,N441,N528);
nand NAND2_150(N576,N444,N531);
nand NAND2_151(N577,N447,N531);
nand NAND2_152(N578,N450,N534);
nand NAND2_153(N579,N453,N534);
nand NAND2_154(N580,N456,N537);
nand NAND2_155(N581,N459,N537);
nand NAND2_156(N582,N462,N540);
nand NAND2_157(N583,N465,N540);
nand NAND2_158(N584,N468,N543);
nand NAND2_159(N585,N471,N543);
nand NAND2_160(N586,N474,N546);
nand NAND2_161(N587,N477,N546);
nand NAND2_162(N588,N480,N549);
nand NAND2_163(N589,N483,N549);
nand NAND2_164(N590,N486,N552);
nand NAND2_165(N591,N489,N552);
nand NAND2_166(N592,N492,N555);
nand NAND2_167(N593,N495,N555);
nand NAND2_168(N594,N498,N558);
nand NAND2_169(N595,N501,N558);
nand NAND2_170(N596,N504,N561);
nand NAND2_171(N597,N507,N561);
nand NAND2_172(N598,N510,N564);
nand NAND2_173(N599,N513,N564);
nand NAND2_174(N600,N516,N567);
nand NAND2_175(N601,N519,N567);
nand NAND2_176(N602,N570,N571);
nand NAND2_177(N607,N572,N573);
nand NAND2_178(N612,N574,N575);
nand NAND2_179(N617,N576,N577);
nand NAND2_180(N622,N578,N579);
nand NAND2_181(N627,N580,N581);
nand NAND2_182(N632,N582,N583);
nand NAND2_183(N637,N584,N585);
nand NAND2_184(N642,N586,N587);
nand NAND2_185(N645,N588,N589);
nand NAND2_186(N648,N590,N591);
nand NAND2_187(N651,N592,N593);
nand NAND2_188(N654,N594,N595);
nand NAND2_189(N657,N596,N597);
nand NAND2_190(N660,N598,N599);
nand NAND2_191(N663,N600,N601);
nand NAND2_192(N666,N602,N607);
nand NAND2_193(N669,N612,N617);
nand NAND2_194(N672,N602,N612);
nand NAND2_195(N675,N607,N617);
nand NAND2_196(N678,N622,N627);
nand NAND2_197(N681,N632,N637);
nand NAND2_198(N684,N622,N632);
nand NAND2_199(N687,N627,N637);
nand NAND2_200(N690,N602,N666);
nand NAND2_201(N691,N607,N666);
nand NAND2_202(N692,N612,N669);
nand NAND2_203(N693,N617,N669);
nand NAND2_204(N694,N602,N672);
nand NAND2_205(N695,N612,N672);
nand NAND2_206(N696,N607,N675);
nand NAND2_207(N697,N617,N675);
nand NAND2_208(N698,N622,N678);
nand NAND2_209(N699,N627,N678);
nand NAND2_210(N700,N632,N681);
nand NAND2_211(N701,N637,N681);
nand NAND2_212(N702,N622,N684);
nand NAND2_213(N703,N632,N684);
nand NAND2_214(N704,N627,N687);
nand NAND2_215(N705,N637,N687);
nand NAND2_216(N706,N690,N691);
nand NAND2_217(N709,N692,N693);
nand NAND2_218(N712,N694,N695);
nand NAND2_219(N715,N696,N697);
nand NAND2_220(N718,N698,N699);
nand NAND2_221(N721,N700,N701);
nand NAND2_222(N724,N702,N703);
nand NAND2_223(N727,N704,N705);
nand NAND2_224(N730,N242,N718);
nand NAND2_225(N733,N245,N721);
nand NAND2_226(N736,N248,N724);
nand NAND2_227(N739,N251,N727);
nand NAND2_228(N742,N254,N706);
nand NAND2_229(N745,N257,N709);
nand NAND2_230(N748,N260,N712);
nand NAND2_231(N751,N263,N715);
nand NAND2_232(N754,N242,N730);
nand NAND2_233(N755,N718,N730);
nand NAND2_234(N756,N245,N733);
nand NAND2_235(N757,N721,N733);
nand NAND2_236(N758,N248,N736);
nand NAND2_237(N759,N724,N736);
nand NAND2_238(N760,N251,N739);
nand NAND2_239(N761,N727,N739);
nand NAND2_240(N762,N254,N742);
nand NAND2_241(N763,N706,N742);
nand NAND2_242(N764,N257,N745);
nand NAND2_243(N765,N709,N745);
nand NAND2_244(N766,N260,N748);
nand NAND2_245(N767,N712,N748);
nand NAND2_246(N768,N263,N751);
nand NAND2_247(N769,N715,N751);
nand NAND2_248(N770,N754,N755);
nand NAND2_249(N773,N756,N757);
nand NAND2_250(N776,N758,N759);
nand NAND2_251(N779,N760,N761);
nand NAND2_252(N782,N762,N763);
nand NAND2_253(N785,N764,N765);
nand NAND2_254(N788,N766,N767);
nand NAND2_255(N791,N768,N769);
nand NAND2_256(N794,N642,N770);
nand NAND2_257(N797,N645,N773);
nand NAND2_258(N800,N648,N776);
nand NAND2_259(N803,N651,N779);
nand NAND2_260(N806,N654,N782);
nand NAND2_261(N809,N657,N785);
nand NAND2_262(N812,N660,N788);
nand NAND2_263(N815,N663,N791);
nand NAND2_264(N818,N642,N794);
nand NAND2_265(N819,N770,N794);
nand NAND2_266(N820,N645,N797);
nand NAND2_267(N821,N773,N797);
nand NAND2_268(N822,N648,N800);
nand NAND2_269(N823,N776,N800);
nand NAND2_270(N824,N651,N803);
nand NAND2_271(N825,N779,N803);
nand NAND2_272(N826,N654,N806);
nand NAND2_273(N827,N782,N806);
nand NAND2_274(N828,N657,N809);
nand NAND2_275(N829,N785,N809);
nand NAND2_276(N830,N660,N812);
nand NAND2_277(N831,N788,N812);
nand NAND2_278(N832,N663,N815);
nand NAND2_279(N833,N791,N815);
nand NAND2_280(N834,N818,N819);
nand NAND2_281(N847,N820,N821);
nand NAND2_282(N860,N822,N823);
nand NAND2_283(N873,N824,N825);
nand NAND2_284(N886,N828,N829);
nand NAND2_285(N899,N832,N833);
nand NAND2_286(N912,N830,N831);
nand NAND2_287(N925,N826,N827);
not NOT1_0(N938,N834);
not NOT1_1(N939,N847);
not NOT1_2(N940,N860);
not NOT1_3(N941,N834);
not NOT1_4(N942,N847);
not NOT1_5(N943,N873);
not NOT1_6(N944,N834);
not NOT1_7(N945,N860);
not NOT1_8(N946,N873);
not NOT1_9(N947,N847);
not NOT1_10(N948,N860);
not NOT1_11(N949,N873);
not NOT1_12(N950,N886);
not NOT1_13(N951,N899);
not NOT1_14(N952,N886);
not NOT1_15(N953,N912);
not NOT1_16(N954,N925);
not NOT1_17(N955,N899);
not NOT1_18(N956,N925);
not NOT1_19(N957,N912);
not NOT1_20(N958,N925);
not NOT1_21(N959,N886);
not NOT1_22(N960,N912);
not NOT1_23(N961,N925);
not NOT1_24(N962,N886);
not NOT1_25(N963,N899);
not NOT1_26(N964,N925);
not NOT1_27(N965,N912);
not NOT1_28(N966,N899);
not NOT1_29(N967,N886);
not NOT1_30(N968,N912);
not NOT1_31(N969,N899);
not NOT1_32(N970,N847);
not NOT1_33(N971,N873);
not NOT1_34(N972,N847);
not NOT1_35(N973,N860);
not NOT1_36(N974,N834);
not NOT1_37(N975,N873);
not NOT1_38(N976,N834);
not NOT1_39(N977,N860);
and AND4_0(N978,N938,N939,N940,N873);
and AND4_1(N979,N941,N942,N860,N943);
and AND4_2(N980,N944,N847,N945,N946);
and AND4_3(N981,N834,N947,N948,N949);
and AND4_4(N982,N958,N959,N960,N899);
and AND4_5(N983,N961,N962,N912,N963);
and AND4_6(N984,N964,N886,N965,N966);
and AND4_7(N985,N925,N967,N968,N969);
or OR4_0(N986,N978,N979,N980,N981);
or OR4_1(N991,N982,N983,N984,N985);
and AND5_0(N996,N925,N950,N912,N951,N986);
and AND5_1(N1001,N925,N952,N953,N899,N986);
and AND5_2(N1006,N954,N886,N912,N955,N986);
and AND5_3(N1011,N956,N886,N957,N899,N986);
and AND5_4(N1016,N834,N970,N860,N971,N991);
and AND5_5(N1021,N834,N972,N973,N873,N991);
and AND5_6(N1026,N974,N847,N860,N975,N991);
and AND5_7(N1031,N976,N847,N977,N873,N991);
and AND2_8(N1036,N834,N996);
and AND2_9(N1039,N847,N996);
and AND2_10(N1042,N860,N996);
and AND2_11(N1045,N873,N996);
and AND2_12(N1048,N834,N1001);
and AND2_13(N1051,N847,N1001);
and AND2_14(N1054,N860,N1001);
and AND2_15(N1057,N873,N1001);
and AND2_16(N1060,N834,N1006);
and AND2_17(N1063,N847,N1006);
and AND2_18(N1066,N860,N1006);
and AND2_19(N1069,N873,N1006);
and AND2_20(N1072,N834,N1011);
and AND2_21(N1075,N847,N1011);
and AND2_22(N1078,N860,N1011);
and AND2_23(N1081,N873,N1011);
and AND2_24(N1084,N925,N1016);
and AND2_25(N1087,N886,N1016);
and AND2_26(N1090,N912,N1016);
and AND2_27(N1093,N899,N1016);
and AND2_28(N1096,N925,N1021);
and AND2_29(N1099,N886,N1021);
and AND2_30(N1102,N912,N1021);
and AND2_31(N1105,N899,N1021);
and AND2_32(N1108,N925,N1026);
and AND2_33(N1111,N886,N1026);
and AND2_34(N1114,N912,N1026);
and AND2_35(N1117,N899,N1026);
and AND2_36(N1120,N925,N1031);
and AND2_37(N1123,N886,N1031);
and AND2_38(N1126,N912,N1031);
and AND2_39(N1129,N899,N1031);
nand NAND2_288(N1132,N1,N1036);
nand NAND2_289(N1135,N8,N1039);
nand NAND2_290(N1138,N15,N1042);
nand NAND2_291(N1141,N22,N1045);
nand NAND2_292(N1144,N29,N1048);
nand NAND2_293(N1147,N36,N1051);
nand NAND2_294(N1150,N43,N1054);
nand NAND2_295(N1153,N50,N1057);
nand NAND2_296(N1156,N57,N1060);
nand NAND2_297(N1159,N64,N1063);
nand NAND2_298(N1162,N71,N1066);
nand NAND2_299(N1165,N78,N1069);
nand NAND2_300(N1168,N85,N1072);
nand NAND2_301(N1171,N92,N1075);
nand NAND2_302(N1174,N99,N1078);
nand NAND2_303(N1177,N106,N1081);
nand NAND2_304(N1180,N113,N1084);
nand NAND2_305(N1183,N120,N1087);
nand NAND2_306(N1186,N127,N1090);
nand NAND2_307(N1189,N134,N1093);
nand NAND2_308(N1192,N141,N1096);
nand NAND2_309(N1195,N148,N1099);
nand NAND2_310(N1198,N155,N1102);
nand NAND2_311(N1201,N162,N1105);
nand NAND2_312(N1204,N169,N1108);
nand NAND2_313(N1207,N176,N1111);
nand NAND2_314(N1210,N183,N1114);
nand NAND2_315(N1213,N190,N1117);
nand NAND2_316(N1216,N197,N1120);
nand NAND2_317(N1219,N204,N1123);
nand NAND2_318(N1222,N211,N1126);
nand NAND2_319(N1225,N218,N1129);
nand NAND2_320(N1228,N1,N1132);
nand NAND2_321(N1229,N1036,N1132);
nand NAND2_322(N1230,N8,N1135);
nand NAND2_323(N1231,N1039,N1135);
nand NAND2_324(N1232,N15,N1138);
nand NAND2_325(N1233,N1042,N1138);
nand NAND2_326(N1234,N22,N1141);
nand NAND2_327(N1235,N1045,N1141);
nand NAND2_328(N1236,N29,N1144);
nand NAND2_329(N1237,N1048,N1144);
nand NAND2_330(N1238,N36,N1147);
nand NAND2_331(N1239,N1051,N1147);
nand NAND2_332(N1240,N43,N1150);
nand NAND2_333(N1241,N1054,N1150);
nand NAND2_334(N1242,N50,N1153);
nand NAND2_335(N1243,N1057,N1153);
nand NAND2_336(N1244,N57,N1156);
nand NAND2_337(N1245,N1060,N1156);
nand NAND2_338(N1246,N64,N1159);
nand NAND2_339(N1247,N1063,N1159);
nand NAND2_340(N1248,N71,N1162);
nand NAND2_341(N1249,N1066,N1162);
nand NAND2_342(N1250,N78,N1165);
nand NAND2_343(N1251,N1069,N1165);
nand NAND2_344(N1252,N85,N1168);
nand NAND2_345(N1253,N1072,N1168);
nand NAND2_346(N1254,N92,N1171);
nand NAND2_347(N1255,N1075,N1171);
nand NAND2_348(N1256,N99,N1174);
nand NAND2_349(N1257,N1078,N1174);
nand NAND2_350(N1258,N106,N1177);
nand NAND2_351(N1259,N1081,N1177);
nand NAND2_352(N1260,N113,N1180);
nand NAND2_353(N1261,N1084,N1180);
nand NAND2_354(N1262,N120,N1183);
nand NAND2_355(N1263,N1087,N1183);
nand NAND2_356(N1264,N127,N1186);
nand NAND2_357(N1265,N1090,N1186);
nand NAND2_358(N1266,N134,N1189);
nand NAND2_359(N1267,N1093,N1189);
nand NAND2_360(N1268,N141,N1192);
nand NAND2_361(N1269,N1096,N1192);
nand NAND2_362(N1270,N148,N1195);
nand NAND2_363(N1271,N1099,N1195);
nand NAND2_364(N1272,N155,N1198);
nand NAND2_365(N1273,N1102,N1198);
nand NAND2_366(N1274,N162,N1201);
nand NAND2_367(N1275,N1105,N1201);
nand NAND2_368(N1276,N169,N1204);
nand NAND2_369(N1277,N1108,N1204);
nand NAND2_370(N1278,N176,N1207);
nand NAND2_371(N1279,N1111,N1207);
nand NAND2_372(N1280,N183,N1210);
nand NAND2_373(N1281,N1114,N1210);
nand NAND2_374(N1282,N190,N1213);
nand NAND2_375(N1283,N1117,N1213);
nand NAND2_376(N1284,N197,N1216);
nand NAND2_377(N1285,N1120,N1216);
nand NAND2_378(N1286,N204,N1219);
nand NAND2_379(N1287,N1123,N1219);
nand NAND2_380(N1288,N211,N1222);
nand NAND2_381(N1289,N1126,N1222);
nand NAND2_382(N1290,N218,N1225);
nand NAND2_383(N1291,N1129,N1225);
nand NAND2_384(N1292,N1228,N1229);
nand NAND2_385(N1293,N1230,N1231);
nand NAND2_386(N1294,N1232,N1233);
nand NAND2_387(N1295,N1234,N1235);
nand NAND2_388(N1296,N1236,N1237);
nand NAND2_389(N1297,N1238,N1239);
nand NAND2_390(N1298,N1240,N1241);
nand NAND2_391(N1299,N1242,N1243);
nand NAND2_392(N1300,N1244,N1245);
nand NAND2_393(N1301,N1246,N1247);
nand NAND2_394(N1302,N1248,N1249);
nand NAND2_395(N1303,N1250,N1251);
nand NAND2_396(N1304,N1252,N1253);
nand NAND2_397(N1305,N1254,N1255);
nand NAND2_398(N1306,N1256,N1257);
nand NAND2_399(N1307,N1258,N1259);
nand NAND2_400(N1308,N1260,N1261);
nand NAND2_401(N1309,N1262,N1263);
nand NAND2_402(N1310,N1264,N1265);
nand NAND2_403(N1311,N1266,N1267);
nand NAND2_404(N1312,N1268,N1269);
nand NAND2_405(N1313,N1270,N1271);
nand NAND2_406(N1314,N1272,N1273);
nand NAND2_407(N1315,N1274,N1275);
nand NAND2_408(N1316,N1276,N1277);
nand NAND2_409(N1317,N1278,N1279);
nand NAND2_410(N1318,N1280,N1281);
nand NAND2_411(N1319,N1282,N1283);
nand NAND2_412(N1320,N1284,N1285);
nand NAND2_413(N1321,N1286,N1287);
nand NAND2_414(N1322,N1288,N1289);
nand NAND2_415(N1323,N1290,N1291);
buf BUFF1_0(N1324,N1292);
buf BUFF1_1(N1325,N1293);
buf BUFF1_2(N1326,N1294);
buf BUFF1_3(N1327,N1295);
buf BUFF1_4(N1328,N1296);
buf BUFF1_5(N1329,N1297);
buf BUFF1_6(N1330,N1298);
buf BUFF1_7(N1331,N1299);
buf BUFF1_8(N1332,N1300);
buf BUFF1_9(N1333,N1301);
buf BUFF1_10(N1334,N1302);
buf BUFF1_11(N1335,N1303);
buf BUFF1_12(N1336,N1304);
buf BUFF1_13(N1337,N1305);
buf BUFF1_14(N1338,N1306);
buf BUFF1_15(N1339,N1307);
buf BUFF1_16(N1340,N1308);
buf BUFF1_17(N1341,N1309);
buf BUFF1_18(N1342,N1310);
buf BUFF1_19(N1343,N1311);
buf BUFF1_20(N1344,N1312);
buf BUFF1_21(N1345,N1313);
buf BUFF1_22(N1346,N1314);
buf BUFF1_23(N1347,N1315);
buf BUFF1_24(N1348,N1316);
buf BUFF1_25(N1349,N1317);
buf BUFF1_26(N1350,N1318);
buf BUFF1_27(N1351,N1319);
buf BUFF1_28(N1352,N1320);
buf BUFF1_29(N1353,N1321);
buf BUFF1_30(N1354,N1322);
buf BUFF1_31(N1355,N1323);

endmodule